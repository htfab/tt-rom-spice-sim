* NGSPICE file created from tt_um_chip_rom.ext - technology: sky130A

.subckt O9_sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt O9_sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt O9_sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt O9_sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt O9_sky130_fd_sc_hd__and4b_1 VGND VPWR VPB VNB C A_N X D B
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o21a_1 VGND VPWR VPB VNB X A1 B1 A2
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__or2_1 VGND VPWR VPB VNB A X B
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__and2b_1 VGND VPWR VPB VNB X A_N B
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__nor2_2 VGND VPWR VPB VNB B Y A
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__buf_2 VPWR VGND VPB VNB X A
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__conb_1 VGND VPWR VPB VNB LO HI
R0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
R1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt O9_sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB A X B C
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__and3_1 VGND VPWR VPB VNB X B A C
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt O9_sky130_fd_sc_hd__a211o_1 VGND VPWR VPB VNB X A2 B1 A1 C1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__nand2_1 VGND VPWR VPB VNB Y B A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o211a_1 VGND VPWR VPB VNB C1 B1 A2 A1 X
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A1 B1 Y A2
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__and2_1 VPWR VGND VPB VNB X B A
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__nor2_1 VGND VPWR VPB VNB B Y A
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB S A1 A0 X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__xnor2_1 VGND VPWR VPB VNB B Y A
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__xor2_1 VPWR VGND VPB VNB B X A
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a31o_1 VGND VPWR VPB VNB A2 B1 A1 A3 X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a311oi_1 VPWR VGND VPB VNB A3 Y C1 B1 A2 A1
X0 Y A1 a_194_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_194_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2 Y C1 a_376_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1725 ps=1.345 w=1 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.112125 ps=0.995 w=0.65 l=0.15
X5 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.115375 ps=1.005 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7 a_376_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.165 ps=1.33 w=1 l=0.15
X8 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a211oi_1 VPWR VGND VPB VNB A1 C1 B1 Y A2
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__clkbuf_4 VGND VPWR VPB VNB X A
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o31a_1 VGND VPWR VPB VNB X A2 B1 A1 A3
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o21ai_1 VGND VPWR VPB VNB A2 A1 B1 Y
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__or3b_1 VGND VPWR VPB VNB A C_N X B
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__or4_1 VPWR VGND VPB VNB C A X B D
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__clkbuf_1 VGND VPWR VPB VNB X A
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__nand2b_1 VGND VPWR VPB VNB Y A_N B
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__clkbuf_2 VGND VPWR VPB VNB A X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a311o_1 VGND VPWR VPB VNB A1 A2 X B1 C1 A3
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.134875 ps=1.065 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.112125 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125125 ps=1.035 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.134875 pd=1.065 as=0.105625 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.1625 ps=1.325 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1425 ps=1.285 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o21ai_2 VGND VPWR VPB VNB B1 Y A2 A1
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__and2b_2 VPWR VGND VPB VNB X B A_N
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.22895 ps=1.745 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22895 pd=1.745 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__buf_1 VGND VPWR VPB VNB X A
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND VPB VNB A X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o21ba_1 VGND VPWR VPB VNB B1_N A1 X A2
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 B2 B1 A1 A2
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__inv_2 VPWR VGND VPB VNB A Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o2bb2a_1 VPWR VGND VPB VNB A1_N X A2_N B2 B1
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o22a_1 VGND VPWR VPB VNB A2 X B1 A1 B2
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a31oi_1 VGND VPWR VPB VNB Y B1 A2 A1 A3
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.118625 ps=1.015 w=0.65 l=0.15
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.06825 ps=0.86 w=0.65 l=0.15
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.105625 ps=0.975 w=0.65 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.1525 ps=1.305 w=1 l=0.15
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o31ai_1 VPWR VGND VPB VNB Y A2 A1 A3 B1
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a221o_1 VPWR VGND VPB VNB X B1 A1 B2 A2 C1
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o221ai_2 VGND VPWR VPB VNB B1 B2 Y A2 A1 C1
X0 Y A2 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_300_47# B2 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 a_300_47# B1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_300_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_734_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7 a_28_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR B1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X11 a_382_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_28_47# B1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_28_47# B2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X15 Y B2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR A1 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_382_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X19 a_734_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB A1 A2 X B2 B1
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a21bo_1 VGND VPWR VPB VNB X A1 B1_N A2
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258375 ps=1.445 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__nor3_1 VGND VPWR VPB VNB C Y A B
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB B X A
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__o221a_1 VGND VPWR VPB VNB A2 X B1 C1 A1 B2
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
.ends

.subckt O9_sky130_fd_sc_hd__a2bb2o_1 VGND VPWR VPB VNB B1 A1_N A2_N X B2
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt tt_um_chip_rom VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_0_27_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_38_81 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_18_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_34_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_200_ VGND VPWR VPWR VGND _023_ _071_ _013_ _078_ net4 O9_sky130_fd_sc_hd__and4b_1
XFILLER_0_33_320 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_131_ VGND VPWR VPWR VGND _051_ net19 _031_ _037_ O9_sky130_fd_sc_hd__o21a_1
XFILLER_0_29_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_191 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_47 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_114_ VGND VPWR VPWR VGND net22 _034_ net27 O9_sky130_fd_sc_hd__or2_1
XFILLER_0_12_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_21_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_34_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_26_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_76 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_37_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_13_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_130_ VGND VPWR VPWR VGND _050_ net20 net21 O9_sky130_fd_sc_hd__and2b_1
XFILLER_0_33_332 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_9_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_63 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_19_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_113_ VGND VPWR VPWR VGND net27 _033_ net22 O9_sky130_fd_sc_hd__nor2_2
XFILLER_0_1_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_21_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_165 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_16_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_50 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_7_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xoutput10 VPWR VGND VPWR VGND uo_out[1] net10 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_27_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_32_249 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_23_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_225__45 VGND VPWR VPWR VGND net45 _225__45/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_37_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_189_ VPWR VGND VPWR VGND net21 _004_ _027_ _047_ O9_sky130_fd_sc_hd__or3_1
XFILLER_0_10_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_19_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_19_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_112_ VGND VPWR VPWR VGND _032_ net25 net22 net27 O9_sky130_fd_sc_hd__and3_1
XFILLER_0_33_130 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_155 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_30_177 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_21_133 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xoutput9 VPWR VGND VPWR VGND uo_out[0] net9 O9_sky130_fd_sc_hd__buf_2
Xoutput11 VPWR VGND VPWR VGND uo_out[2] net11 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_23_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_13_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_24_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_188_ VGND VPWR VPWR VGND _003_ _000_ _001_ net16 _002_ O9_sky130_fd_sc_hd__a211o_1
XFILLER_0_34_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_142 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_111_ VGND VPWR VPWR VGND _031_ net27 net25 O9_sky130_fd_sc_hd__nand2_1
XFILLER_0_8_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_131 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_24_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_145 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_178 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_32_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_204 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xoutput12 VPWR VGND VPWR VGND uo_out[3] net12 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_7_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_26_204 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_17_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_38_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_36_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_216__36 VGND VPWR VPWR VGND net36 _216__36/HI O9_sky130_fd_sc_hd__conb_1
X_187_ VGND VPWR VPWR VGND _025_ net20 _033_ _032_ _002_ O9_sky130_fd_sc_hd__o211a_1
X_110_ VPWR VGND VPWR VGND net25 net18 _030_ _029_ O9_sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_176 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_154 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_67 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_24_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_21_157 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_16_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_32_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_216 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
Xoutput13 VPWR VGND VPWR VGND uo_out[4] net13 O9_sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_17_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_54 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_39 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_24_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_10_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_186_ VPWR VGND VPWR VGND _001_ _054_ _025_ O9_sky130_fd_sc_hd__and2_1
XFILLER_0_18_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_188 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_42 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_24_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_169_ VGND VPWR VPWR VGND _085_ _086_ _084_ O9_sky130_fd_sc_hd__nor2_1
XFILLER_0_38_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_18_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xoutput14 VPWR VGND VPWR VGND uo_out[5] net14 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_1_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_71 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_1_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_18_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_5_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_185_ VGND VPWR VPWR VGND _099_ _100_ net17 _000_ O9_sky130_fd_sc_hd__mux2_1
XFILLER_0_2_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_318 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_221__41 VGND VPWR VPWR VGND net41 _221__41/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_18_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_21_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_168_ VGND VPWR VPWR VGND net23 _024_ _028_ _085_ O9_sky130_fd_sc_hd__mux2_1
XFILLER_0_38_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xoutput15 VPWR VGND VPWR VGND uo_out[6] net15 O9_sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_229 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_25_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_25_295 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_30_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_11 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_1_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_36_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_184_ VGND VPWR VPWR VGND _100_ net24 _023_ _047_ O9_sky130_fd_sc_hd__o21a_1
XFILLER_0_19_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_167_ VPWR VGND VPWR VGND net21 net20 _084_ _083_ O9_sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_249 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_21_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_29_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_219_ VPWR VGND VPWR VGND uio_out[2] net39 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_29_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_171 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_241 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_19_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_1_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_58 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_9_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_193 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_36_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_183_ VGND VPWR VPWR VGND _083_ _099_ _057_ O9_sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_18_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_212__32 VGND VPWR VPWR VGND net32 _212__32/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_21_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_114 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_166_ VPWR VGND VPWR VGND net28 _083_ net26 O9_sky130_fd_sc_hd__xor2_1
XFILLER_0_1_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_46 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_16_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_218_ VPWR VGND VPWR VGND uio_out[1] net38 O9_sky130_fd_sc_hd__buf_2
X_149_ VGND VPWR VPWR VGND _031_ net17 net24 _039_ _068_ O9_sky130_fd_sc_hd__a31o_1
XFILLER_0_20_183 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_34_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_212 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_245 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_289 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_9_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Left_75 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_59 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_24_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_307 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_182_ VPWR VGND VPWR VGND _091_ net12 net8 _098_ _090_ _026_ O9_sky130_fd_sc_hd__a311oi_1
XFILLER_0_36_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_19_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_27_134 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_18_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_165_ VPWR VGND VPWR VGND net6 _082_ _077_ net11 _075_ O9_sky130_fd_sc_hd__a211oi_1
XFILLER_0_21_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_62 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_11_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_118 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_37_262 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_217_ VPWR VGND VPWR VGND uio_out[0] net37 O9_sky130_fd_sc_hd__buf_2
X_148_ VPWR VGND VPWR VGND _031_ net24 _045_ _067_ _039_ O9_sky130_fd_sc_hd__a211oi_1
XFILLER_0_34_287 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_27_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_17_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_257 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_13_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_224 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_25 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_219__39 VGND VPWR VPWR VGND net39 _219__39/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_27_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xfanout20 VGND VPWR VPWR VGND net20 net4 O9_sky130_fd_sc_hd__clkbuf_4
X_181_ VGND VPWR VPWR VGND _098_ _094_ net7 net6 _097_ O9_sky130_fd_sc_hd__o31a_1
XFILLER_0_10_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_146 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_21_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_164_ VGND VPWR VPWR VGND _082_ _079_ net7 _081_ O9_sky130_fd_sc_hd__and3_1
XFILLER_0_1_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_15_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_37_285 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_216_ VPWR VGND VPWR VGND uio_oe[7] net36 O9_sky130_fd_sc_hd__buf_2
X_147_ VGND VPWR VPWR VGND _065_ _029_ _026_ _066_ O9_sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_141 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_299 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_27_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_3_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_22_236 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xfanout21 VPWR VGND VPWR VGND net21 net24 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_36_114 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_180_ VGND VPWR VPWR VGND _097_ _095_ net18 _096_ O9_sky130_fd_sc_hd__o21a_1
XFILLER_0_24_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_158 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_27_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_163_ VGND VPWR VPWR VGND _023_ _080_ _081_ _049_ O9_sky130_fd_sc_hd__or3b_1
XFILLER_0_1_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_23_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_38_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_37_297 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_37_220 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
X_215_ VPWR VGND VPWR VGND uio_oe[6] net35 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_4_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_146_ VPWR VGND VPWR VGND _040_ net17 _065_ net16 _045_ O9_sky130_fd_sc_hd__or4_1
XFILLER_0_12_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_7_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_129_ VGND VPWR VPWR VGND _046_ _049_ _037_ O9_sky130_fd_sc_hd__nor2_1
XFILLER_0_33_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_248 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_13_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_224__44 VGND VPWR VPWR VGND net44 _224__44/HI O9_sky130_fd_sc_hd__conb_1
Xfanout22 VPWR VGND VPWR VGND net22 net24 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_3_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_162_ VGND VPWR VPWR VGND net27 net22 net19 _080_ O9_sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
Xinput1 VGND VPWR VPWR VGND net1 ui_in[0] O9_sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_214_ VPWR VGND VPWR VGND uio_oe[5] net34 O9_sky130_fd_sc_hd__buf_2
X_145_ VGND VPWR VPWR VGND _064_ _061_ net16 _063_ O9_sky130_fd_sc_hd__o21a_1
XFILLER_0_20_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_66 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_7_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_210 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_128_ VGND VPWR VPWR VGND _048_ net26 net28 O9_sky130_fd_sc_hd__nand2b_1
XFILLER_0_17_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_38_17 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_13_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_53 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_8_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xfanout23 VGND VPWR VPWR VGND net24 net23 O9_sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_35_193 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_25_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_1_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_161_ VGND VPWR VPWR VGND _022_ _034_ _079_ _059_ net18 _078_ O9_sky130_fd_sc_hd__a311o_1
XFILLER_0_17_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xinput2 VGND VPWR VPWR VGND net2 ui_in[1] O9_sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_37_277 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_213_ VPWR VGND VPWR VGND uio_oe[4] net33 O9_sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_2_Left_41 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_144_ VGND VPWR VPWR VGND _039_ _034_ _062_ _063_ O9_sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_22_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_222 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_127_ VGND VPWR VPWR VGND _047_ net25 net27 O9_sky130_fd_sc_hd__and2b_1
XFILLER_0_33_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_38_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_8_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_70 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_14_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_191 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_5_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_320 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xfanout24 VGND VPWR VPWR VGND net3 net24 O9_sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_128 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_215__35 VGND VPWR VPWR VGND net35 _215__35/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_35_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_23_301 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_5_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_17_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_160_ VGND VPWR VPWR VGND net23 _078_ net27 net25 O9_sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
Xinput3 VGND VPWR VPWR VGND net3 ui_in[2] O9_sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_14_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_212_ VPWR VGND VPWR VGND uio_oe[3] net32 O9_sky130_fd_sc_hd__buf_2
X_143_ VPWR VGND VPWR VGND _040_ net18 _062_ _033_ _057_ O9_sky130_fd_sc_hd__or4_1
XFILLER_0_22_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_234 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_126_ VGND VPWR VPWR VGND net27 _046_ net25 O9_sky130_fd_sc_hd__nor2_2
XFILLER_0_24_292 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_218 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_109_ VPWR VGND VPWR VGND _029_ net21 net28 O9_sky130_fd_sc_hd__and2b_2
XFILLER_0_28_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_8_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_332 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_5_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xfanout25 VPWR VGND VPWR VGND net25 net26 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_29_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_313 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_32_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xinput4 VGND VPWR VPWR VGND net4 ui_in[3] O9_sky130_fd_sc_hd__buf_1
XFILLER_0_36_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_211_ VPWR VGND VPWR VGND uio_oe[2] net31 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_9_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_142_ VGND VPWR VPWR VGND net18 _060_ _059_ _046_ _061_ O9_sky130_fd_sc_hd__o211a_1
XFILLER_0_22_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_246 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_11_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_249 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_125_ VGND VPWR VPWR VGND _024_ _045_ net19 O9_sky130_fd_sc_hd__nor2_2
XFILLER_0_25_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_24_260 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_241 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_108_ VGND VPWR VPWR VGND _028_ net27 net25 O9_sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_5_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_57 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_30_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xfanout26 VGND VPWR VPWR VGND net26 net2 O9_sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_160 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_29_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_325 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_26_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_220__40 VGND VPWR VPWR VGND net40 _220__40/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_32_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_32_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xinput5 VGND VPWR VPWR VGND net5 ui_in[4] O9_sky130_fd_sc_hd__buf_1
XFILLER_0_36_97 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_36_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
X_210_ VPWR VGND VPWR VGND uio_oe[1] net30 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_9_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_141_ VGND VPWR VPWR VGND _060_ _046_ net19 O9_sky130_fd_sc_hd__nand2_1
XFILLER_0_22_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_45 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_124_ VGND VPWR VPWR VGND _043_ net7 net16 _044_ O9_sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_206 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_272 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_107_ VGND VPWR VPWR VGND _027_ net28 net26 O9_sky130_fd_sc_hd__and2b_1
XFILLER_0_0_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_331 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_8_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_183 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_5_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_30_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
Xfanout16 VGND VPWR VPWR VGND net16 net6 O9_sky130_fd_sc_hd__clkbuf_4
Xfanout27 VGND VPWR VPWR VGND net27 net28 O9_sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_35_Left_74 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_11_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
Xinput6 VPWR VGND VPWR VGND ui_in[5] net6 O9_sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_36_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_21 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_6_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_14_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_140_ VGND VPWR VPWR VGND _057_ net22 _059_ _027_ O9_sky130_fd_sc_hd__o21ba_1
XFILLER_0_20_159 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_11_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_61 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_123_ VGND VPWR VPWR VGND _043_ _042_ _030_ _035_ net18 _024_ O9_sky130_fd_sc_hd__a32o_1
XFILLER_0_25_218 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_24_284 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_28_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_106_ VPWR VGND VPWR VGND net7 _026_ O9_sky130_fd_sc_hd__inv_2
XFILLER_0_0_137 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_28_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_8_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_302 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_151 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
Xfanout17 VPWR VGND VPWR VGND net17 net5 O9_sky130_fd_sc_hd__buf_2
Xfanout28 VPWR VGND VPWR VGND net28 net1 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_32_327 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_26_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_211__31 VGND VPWR VPWR VGND net31 _211__31/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_11_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_11 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
Xinput7 VPWR VGND VPWR VGND net7 ui_in[6] O9_sky130_fd_sc_hd__buf_2
XFILLER_0_36_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_37_249 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_20_149 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_199_ VPWR VGND VPWR VGND _026_ net8 _012_ net14 _010_ O9_sky130_fd_sc_hd__a211oi_1
XFILLER_0_36_282 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_260 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_122_ VPWR VGND VPWR VGND net19 _042_ _037_ net23 _039_ O9_sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_17_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_30_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_105_ VPWR VGND VPWR VGND net16 _025_ O9_sky130_fd_sc_hd__inv_2
XFILLER_0_21_266 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xfanout18 VPWR VGND VPWR VGND net18 net5 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_29_152 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_25_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xinput8 VGND VPWR VPWR VGND ui_in[7] net8 O9_sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_294 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_198_ VGND VPWR VPWR VGND _012_ net16 net7 _011_ O9_sky130_fd_sc_hd__o21a_1
XFILLER_0_19_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_34_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_27_272 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_121_ VGND VPWR VPWR VGND net22 _041_ net26 O9_sky130_fd_sc_hd__or2_1
XFILLER_0_0_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_30_289 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_104_ VPWR VGND VPWR VGND net27 _024_ O9_sky130_fd_sc_hd__inv_2
XFILLER_0_12_245 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_12_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_218__38 VGND VPWR VPWR VGND net38 _218__38/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_38_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_175 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
Xfanout19 VGND VPWR VPWR VGND net19 net20 O9_sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_120 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_197_ VGND VPWR VPWR VGND net20 net21 _046_ net17 _011_ O9_sky130_fd_sc_hd__o211a_1
XFILLER_0_3_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_120_ VGND VPWR VPWR VGND net26 _040_ net21 O9_sky130_fd_sc_hd__nor2_1
XFILLER_0_17_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_65 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_33_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_49 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_24_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_302 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_21_202 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_103_ VPWR VGND VPWR VGND net17 _023_ O9_sky130_fd_sc_hd__inv_2
XFILLER_0_26_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_30_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_29_132 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_52 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_23_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_37_208 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_241 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_196_ VGND VPWR VPWR VGND _088_ _001_ net16 _009_ _010_ O9_sky130_fd_sc_hd__a31o_1
XFILLER_0_2_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_200 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_40 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_17_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_179_ VGND VPWR VPWR VGND _038_ _096_ _041_ _033_ net4 O9_sky130_fd_sc_hd__o22a_1
XFILLER_0_3_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_102_ VPWR VGND VPWR VGND net19 _022_ O9_sky130_fd_sc_hd__inv_2
XFILLER_0_28_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_209__29 VGND VPWR VPWR VGND net29 _209__29/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_17_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_144 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_4_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
X_223__43 VGND VPWR VPWR VGND net43 _223__43/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_35_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_136 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_5_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_10_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_13_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_195_ VPWR VGND VPWR VGND _027_ _022_ _023_ _009_ O9_sky130_fd_sc_hd__a21o_1
XFILLER_0_27_231 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_212 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_178_ VGND VPWR VPWR VGND _078_ _095_ _022_ O9_sky130_fd_sc_hd__nor2_1
XFILLER_0_23_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_326 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_101_ VPWR VGND VPWR VGND net8 _021_ O9_sky130_fd_sc_hd__inv_2
XFILLER_0_0_109 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_4_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_29_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_210 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_194_ VPWR VGND VPWR VGND _026_ net8 _008_ net13 _003_ O9_sky130_fd_sc_hd__a211oi_1
XFILLER_0_2_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_243 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_177_ VGND VPWR VPWR VGND _094_ _055_ _093_ _092_ O9_sky130_fd_sc_hd__o21a_1
XFILLER_0_30_249 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_3_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_11_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_35_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_214__34 VGND VPWR VPWR VGND net34 _214__34/HI O9_sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_26_Right_26 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_34_193 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_300 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_5_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_56 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_182 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_9_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_222 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_193_ VGND VPWR VPWR VGND _008_ _026_ _005_ _025_ _007_ O9_sky130_fd_sc_hd__a31oi_1
XFILLER_0_2_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_176_ VGND VPWR VPWR VGND _093_ _047_ _080_ net22 _037_ O9_sky130_fd_sc_hd__a211o_1
XFILLER_0_15_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_44 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_28_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_159_ VPWR VGND VPWR VGND _077_ net7 net6 _076_ _056_ O9_sky130_fd_sc_hd__o31ai_1
XFILLER_0_11_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_320 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_117 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_1_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_9_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_194 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_32_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_73 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_6_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_192_ VGND VPWR VPWR VGND _006_ _058_ net17 _007_ O9_sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_33_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_175_ VGND VPWR VPWR VGND _092_ _023_ net22 _028_ O9_sky130_fd_sc_hd__and3_1
XFILLER_0_15_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_60 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_21_218 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_8_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_158_ VGND VPWR VPWR VGND _076_ _028_ _033_ net22 _037_ O9_sky130_fd_sc_hd__a211o_1
XFILLER_0_18_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_38_159 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_38_137 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_34_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_332 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_20_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_313 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_22_165 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_26_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_191_ VGND VPWR VPWR VGND _039_ _006_ _029_ O9_sky130_fd_sc_hd__nor2_1
XFILLER_0_12_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_174_ VGND VPWR VPWR VGND _091_ _029_ _054_ net26 net16 O9_sky130_fd_sc_hd__a211o_1
XFILLER_0_2_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_29_319 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_157_ VPWR VGND VPWR VGND _075_ _074_ net18 _030_ _073_ net7 O9_sky130_fd_sc_hd__a221o_1
XFILLER_0_18_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_209_ VPWR VGND VPWR VGND uio_oe[0] net29 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_20_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_3_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_25_130 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_22_188 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_9_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_190_ VPWR VGND VPWR VGND _005_ _084_ _036_ _004_ _048_ net17 O9_sky130_fd_sc_hd__a221o_1
XFILLER_0_12_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_27_203 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_291 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_173_ VGND VPWR VPWR VGND _088_ _089_ _090_ _087_ _086_ net16 O9_sky130_fd_sc_hd__o221ai_2
XFILLER_0_32_283 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_225_ VPWR VGND VPWR VGND uo_out[7] net45 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_12_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_156_ VPWR VGND VPWR VGND _040_ _022_ _058_ _074_ O9_sky130_fd_sc_hd__a21o_1
XFILLER_0_20_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_48 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_37_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_139_ VGND VPWR VPWR VGND _058_ net21 net20 _027_ O9_sky130_fd_sc_hd__o21a_1
X_208_ VPWR VGND VPWR VGND _026_ net8 _015_ net15 _020_ O9_sky130_fd_sc_hd__a211oi_1
XFILLER_0_16_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_3_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_34_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_142 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_0_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_210__30 VGND VPWR VPWR VGND net30 _210__30/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_26_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_215 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_35_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_172_ VGND VPWR VPWR VGND _089_ _037_ _045_ O9_sky130_fd_sc_hd__and2b_1
XFILLER_0_32_295 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_224_ VPWR VGND VPWR VGND uio_out[7] net44 O9_sky130_fd_sc_hd__buf_2
X_155_ VPWR VGND VPWR VGND _041_ _045_ _073_ net19 _072_ O9_sky130_fd_sc_hd__a22o_1
XFILLER_0_18_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_64 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_34_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_207_ VGND VPWR VPWR VGND _025_ _019_ _018_ _020_ O9_sky130_fd_sc_hd__mux2_1
X_138_ VGND VPWR VPWR VGND _057_ net21 net20 net26 O9_sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_305 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_3_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_34_121 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_34_132 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_13_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_51 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_16_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_26_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_13_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_190 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_249 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_35_293 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_26_271 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_171_ VGND VPWR VPWR VGND net20 net17 net21 _046_ _088_ O9_sky130_fd_sc_hd__a31o_1
XFILLER_0_32_241 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_223_ VPWR VGND VPWR VGND uio_out[6] net43 O9_sky130_fd_sc_hd__buf_2
X_154_ VGND VPWR VPWR VGND _032_ _072_ _071_ O9_sky130_fd_sc_hd__or2_1
XFILLER_0_20_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_7_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_3 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_217__37 VGND VPWR VPWR VGND net37 _217__37/HI O9_sky130_fd_sc_hd__conb_1
X_137_ VGND VPWR VPWR VGND _044_ _056_ _053_ _026_ net9 O9_sky130_fd_sc_hd__o211a_1
XFILLER_0_37_196 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_206_ VPWR VGND VPWR VGND _019_ _036_ _022_ _047_ _027_ _054_ O9_sky130_fd_sc_hd__a221o_1
XFILLER_0_28_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_16_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_16_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_283 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_24_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_170_ VPWR VGND VPWR VGND _085_ _084_ _023_ _087_ O9_sky130_fd_sc_hd__a21o_1
XFILLER_0_17_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_231 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_222_ VPWR VGND VPWR VGND uio_out[5] net42 O9_sky130_fd_sc_hd__buf_2
X_153_ VGND VPWR VPWR VGND net28 _071_ net23 net26 O9_sky130_fd_sc_hd__nor3_1
XFILLER_0_20_212 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_28_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_38_109 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_29_109 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_136_ VGND VPWR VPWR VGND _056_ net7 _021_ net16 _055_ O9_sky130_fd_sc_hd__o31a_1
XFILLER_0_4_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_205_ VPWR VGND VPWR VGND net17 _018_ _016_ _088_ _017_ O9_sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_34_156 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
X_119_ VPWR VGND VPWR VGND net19 _039_ net25 O9_sky130_fd_sc_hd__or2_2
XFILLER_0_8_301 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_16_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_192 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_13_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_12_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_17_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_221_ VPWR VGND VPWR VGND uio_out[4] net41 O9_sky130_fd_sc_hd__buf_2
X_152_ VGND VPWR VPWR VGND _066_ net10 _070_ _021_ _064_ _026_ O9_sky130_fd_sc_hd__o221a_1
XFILLER_0_9_281 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_224 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_204_ VGND VPWR VPWR VGND _017_ _050_ net20 _037_ net26 net28 O9_sky130_fd_sc_hd__a32o_1
XFILLER_0_20_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_68 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_135_ VGND VPWR VPWR VGND _055_ net19 _023_ _037_ O9_sky130_fd_sc_hd__o21a_1
XFILLER_0_29_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_222__42 VGND VPWR VPWR VGND net42 _222__42/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_30_330 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_15_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_118_ VGND VPWR VPWR VGND net19 _038_ net25 O9_sky130_fd_sc_hd__nor2_1
XFILLER_0_31_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_31_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_38_271 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_5_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_55 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_8_165 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_241 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_32_211 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_266 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_220_ VPWR VGND VPWR VGND uio_out[3] net40 O9_sky130_fd_sc_hd__buf_2
XFILLER_0_9_293 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_151_ VGND VPWR VPWR VGND _068_ _070_ _069_ _025_ _067_ _023_ O9_sky130_fd_sc_hd__o221a_1
XFILLER_0_18_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_236 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_43 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
X_203_ VPWR VGND VPWR VGND _036_ _016_ _048_ _050_ O9_sky130_fd_sc_hd__or3_1
X_134_ VGND VPWR VPWR VGND net17 _054_ _050_ O9_sky130_fd_sc_hd__or2_1
XFILLER_0_29_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_34_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_69 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_15_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_117_ VPWR VGND VPWR VGND _037_ net25 net22 O9_sky130_fd_sc_hd__and2b_2
XFILLER_0_25_169 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_31_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_2_309 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_72 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_10_109 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_220 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_5_169 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_26_297 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_32_223 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_23_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_245 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_23_256 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_3_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_1_161 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_150_ VGND VPWR VPWR VGND _050_ net28 _057_ _069_ _047_ O9_sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_20_248 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_16_Right_16 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_11_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Right_34 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_25_307 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
X_133_ VGND VPWR VPWR VGND _053_ _045_ _052_ net18 _049_ O9_sky130_fd_sc_hd__o31a_1
X_202_ VGND VPWR VPWR VGND _015_ _013_ net7 net6 _014_ O9_sky130_fd_sc_hd__o31a_1
XFILLER_0_29_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_19_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_213__33 VGND VPWR VPWR VGND net33 _213__33/HI O9_sky130_fd_sc_hd__conb_1
XFILLER_0_15_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_116_ VGND VPWR VPWR VGND _036_ net21 net20 O9_sky130_fd_sc_hd__and2b_1
XFILLER_0_25_159 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_31_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_6_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_12_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_27_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_0_3 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_37_124 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_37_179 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_132_ VGND VPWR VPWR VGND _051_ _032_ net18 _052_ O9_sky130_fd_sc_hd__o21ai_1
X_201_ VGND VPWR VPWR VGND _028_ _014_ _029_ net18 net23 _039_ O9_sky130_fd_sc_hd__o221a_1
XFILLER_0_29_27 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_300 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_25_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
X_115_ VGND VPWR VPWR VGND _033_ _032_ _022_ _035_ O9_sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_249 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_3
XFILLER_0_1_93 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_30_130 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_8
XFILLER_0_38_263 VGND VPWR VPWR VGND O9_sky130_fd_sc_hd__decap_4
XFILLER_0_29_274 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
XFILLER_0_12_141 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VPWR VPWR VGND O9_sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VPWR VGND VPWR VGND O9_sky130_fd_sc_hd__decap_6
.ends


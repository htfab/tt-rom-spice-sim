* Extracted by KLayout with SG13G2 LVS runset on : 11/11/2024 01:28

.SUBCKT tt_um_chip_rom VGND VPWR ui_in[4] ui_in[0] ui_in[3] ui_in[2] ui_in[1]
+ ui_in[5] ui_in[6] ui_in[7] uo_out[2] uo_out[4] uo_out[0] uo_out[7] uo_out[6]
+ uo_out[3] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2]
+ uio_oe[1] uio_oe[0] uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3]
+ uio_out[2] uio_out[1] uio_out[0] uo_out[5] uo_out[1]
X$7 VGND VPWR sg13g2_decap_8
X$8 VGND VPWR sg13g2_decap_8
X$9 VGND VPWR sg13g2_decap_8
X$10 VGND VPWR sg13g2_decap_8
X$11 VGND VPWR sg13g2_decap_8
X$12 VGND VPWR sg13g2_decap_8
X$14 VGND VPWR sg13g2_decap_8
X$15 VGND VPWR sg13g2_decap_8
X$16 VGND VPWR sg13g2_decap_8
X$17 VGND VPWR sg13g2_decap_8
X$18 VGND VPWR sg13g2_decap_8
X$19 VGND VPWR sg13g2_decap_8
X$20 VGND VPWR sg13g2_decap_8
X$21 VGND VPWR sg13g2_decap_8
X$22 VGND VPWR sg13g2_decap_8
X$23 VGND VPWR sg13g2_decap_8
X$24 VGND VPWR sg13g2_decap_8
X$25 VGND VPWR sg13g2_decap_8
X$26 VGND VPWR sg13g2_decap_8
X$27 VGND VPWR sg13g2_decap_8
X$28 VGND VPWR sg13g2_decap_8
X$29 VGND VPWR sg13g2_decap_8
X$30 VGND VPWR sg13g2_decap_8
X$31 VGND VPWR sg13g2_decap_8
X$32 VGND VPWR sg13g2_decap_8
X$33 VGND VPWR sg13g2_decap_8
X$34 VGND VPWR sg13g2_decap_8
X$35 VGND VPWR sg13g2_decap_8
X$36 VGND VPWR sg13g2_decap_8
X$38 VGND VPWR sg13g2_decap_8
X$39 VGND VPWR sg13g2_decap_8
X$40 VGND VPWR sg13g2_decap_8
X$41 VGND VPWR sg13g2_decap_8
X$42 VGND VPWR sg13g2_decap_8
X$43 VGND VPWR sg13g2_decap_8
X$44 VGND VPWR sg13g2_decap_8
X$45 VGND VPWR sg13g2_decap_8
X$46 VGND VPWR sg13g2_decap_8
X$47 VGND VPWR sg13g2_decap_8
X$48 VGND VPWR sg13g2_decap_8
X$49 VGND VPWR sg13g2_decap_8
X$50 VGND VPWR sg13g2_decap_8
X$51 VGND VPWR sg13g2_decap_8
X$52 VGND VPWR sg13g2_decap_8
X$53 VGND VPWR sg13g2_decap_8
X$54 VGND VPWR sg13g2_decap_8
X$55 VGND VPWR sg13g2_decap_8
X$56 VGND VPWR sg13g2_decap_8
X$57 VGND VPWR sg13g2_decap_8
X$58 VGND VPWR sg13g2_decap_8
X$59 VGND VPWR sg13g2_decap_8
X$61 VGND VPWR sg13g2_decap_8
X$62 VGND VPWR sg13g2_decap_8
X$63 VGND VPWR sg13g2_decap_8
X$64 VGND VPWR sg13g2_decap_8
X$65 VGND VPWR sg13g2_decap_8
X$66 VGND VPWR sg13g2_decap_8
X$67 VGND VPWR sg13g2_decap_8
X$68 VGND VPWR sg13g2_decap_8
X$69 VGND VPWR sg13g2_decap_8
X$70 VGND VPWR sg13g2_decap_8
X$73 VGND VPWR sg13g2_decap_8
X$74 VGND VPWR sg13g2_decap_8
X$75 VGND VPWR sg13g2_decap_8
X$76 VGND VPWR sg13g2_decap_8
X$77 VGND VPWR sg13g2_decap_8
X$78 VGND VPWR sg13g2_decap_8
X$82 VGND VPWR sg13g2_decap_8
X$83 VGND VPWR sg13g2_decap_8
X$84 VGND VPWR sg13g2_decap_8
X$85 VGND VPWR sg13g2_decap_8
X$86 VGND VPWR sg13g2_decap_8
X$87 VGND VPWR sg13g2_decap_8
X$88 VGND VPWR sg13g2_decap_8
X$89 VGND VPWR sg13g2_decap_8
X$90 VGND VPWR sg13g2_decap_8
X$91 VGND VPWR sg13g2_decap_8
X$92 VGND VPWR sg13g2_decap_8
X$93 VGND VPWR sg13g2_decap_8
X$94 VGND VPWR sg13g2_decap_8
X$95 VGND VPWR sg13g2_decap_8
X$96 VGND VPWR sg13g2_decap_8
X$97 VGND VPWR sg13g2_decap_8
X$98 VGND VPWR sg13g2_decap_8
X$99 VGND VPWR sg13g2_decap_8
X$100 VGND VPWR sg13g2_decap_8
X$101 VGND VPWR sg13g2_decap_8
X$102 VGND VPWR sg13g2_decap_8
X$103 VGND VPWR sg13g2_decap_8
X$104 VGND VPWR sg13g2_decap_8
X$108 VGND VPWR sg13g2_decap_8
X$109 VGND VPWR sg13g2_decap_8
X$110 VGND VPWR sg13g2_decap_8
X$111 VGND VPWR sg13g2_decap_8
X$112 VGND VPWR sg13g2_decap_8
X$113 VGND VPWR sg13g2_decap_8
X$114 VGND VPWR sg13g2_decap_8
X$115 VGND VPWR sg13g2_decap_8
X$116 VGND VPWR sg13g2_decap_8
X$117 VGND VPWR sg13g2_decap_8
X$118 VGND VPWR sg13g2_decap_8
X$119 VGND VPWR sg13g2_decap_8
X$120 VGND VPWR sg13g2_decap_8
X$121 VGND VPWR sg13g2_decap_8
X$122 VGND VPWR sg13g2_decap_8
X$123 VGND VPWR sg13g2_decap_8
X$124 VGND VPWR sg13g2_decap_8
X$125 VGND VPWR sg13g2_decap_8
X$126 VGND VPWR sg13g2_decap_8
X$127 VGND VPWR sg13g2_decap_8
X$128 VGND VPWR sg13g2_decap_8
X$129 VGND VPWR sg13g2_decap_8
X$133 VGND VPWR sg13g2_decap_8
X$134 VGND VPWR sg13g2_decap_8
X$135 VGND VPWR sg13g2_decap_8
X$136 VGND VPWR sg13g2_decap_8
X$137 VGND VPWR sg13g2_decap_8
X$138 VGND VPWR sg13g2_decap_8
X$139 VGND VPWR sg13g2_decap_8
X$140 VGND VPWR sg13g2_decap_8
X$141 VGND VPWR sg13g2_decap_8
X$142 VGND VPWR sg13g2_decap_8
X$145 VGND VPWR sg13g2_decap_8
X$146 VGND VPWR sg13g2_decap_8
X$147 VGND VPWR sg13g2_decap_8
X$148 VGND VPWR sg13g2_decap_8
X$149 VGND VPWR sg13g2_decap_8
X$150 VGND VPWR sg13g2_decap_8
X$151 VGND VPWR sg13g2_decap_8
X$152 VGND VPWR sg13g2_decap_8
X$157 VGND VPWR sg13g2_decap_8
X$158 VGND VPWR sg13g2_decap_8
X$159 VGND VPWR sg13g2_decap_8
X$160 VGND VPWR sg13g2_decap_8
X$165 VGND VPWR sg13g2_decap_8
X$166 VGND VPWR sg13g2_decap_8
X$167 VGND VPWR sg13g2_decap_8
X$168 VGND VPWR sg13g2_decap_8
X$169 VGND VPWR sg13g2_decap_8
X$170 VGND VPWR sg13g2_decap_8
X$171 VGND VPWR sg13g2_decap_8
X$172 VGND VPWR sg13g2_decap_8
X$173 VGND VPWR sg13g2_decap_8
X$174 VGND VPWR sg13g2_decap_8
X$175 VGND VPWR sg13g2_decap_8
X$176 VGND VPWR sg13g2_decap_8
X$177 VGND VPWR sg13g2_decap_8
X$178 VGND VPWR sg13g2_decap_8
X$179 VGND VPWR sg13g2_decap_8
X$180 VGND VPWR sg13g2_decap_8
X$181 VGND VPWR sg13g2_decap_8
X$182 VGND VPWR sg13g2_decap_8
X$183 VGND VPWR sg13g2_decap_8
X$184 VGND VPWR sg13g2_decap_8
X$185 VGND VPWR sg13g2_decap_8
X$186 VGND VPWR sg13g2_decap_8
X$187 VGND VPWR sg13g2_decap_8
X$188 VGND VPWR sg13g2_decap_8
X$189 VGND VPWR sg13g2_decap_8
X$190 VGND VPWR sg13g2_decap_8
X$191 VGND VPWR sg13g2_decap_8
X$192 VGND VPWR sg13g2_decap_8
X$193 VGND VPWR sg13g2_decap_8
X$194 VGND VPWR sg13g2_decap_8
X$195 VGND VPWR sg13g2_decap_8
X$196 VGND VPWR sg13g2_decap_8
X$197 VGND VPWR sg13g2_decap_8
X$198 VGND VPWR sg13g2_decap_8
X$199 VGND VPWR sg13g2_decap_8
X$200 VGND VPWR sg13g2_decap_8
X$201 VGND VPWR sg13g2_decap_8
X$202 VGND VPWR sg13g2_decap_8
X$203 VGND VPWR sg13g2_decap_8
X$204 VGND VPWR sg13g2_decap_8
X$205 VGND VPWR sg13g2_decap_8
X$206 VGND VPWR sg13g2_decap_8
X$211 VGND VPWR sg13g2_decap_8
X$212 VGND VPWR sg13g2_decap_8
X$213 VGND VPWR sg13g2_decap_8
X$214 VGND VPWR sg13g2_decap_8
X$219 VGND VPWR sg13g2_decap_8
X$220 VGND VPWR sg13g2_decap_8
X$221 VGND VPWR sg13g2_decap_8
X$222 VGND VPWR sg13g2_decap_8
X$223 VGND VPWR sg13g2_decap_8
X$224 VGND VPWR sg13g2_decap_8
X$225 VGND VPWR sg13g2_decap_8
X$226 VGND VPWR sg13g2_decap_8
X$227 VGND VPWR sg13g2_decap_8
X$228 VGND VPWR sg13g2_decap_8
X$229 VGND VPWR sg13g2_decap_8
X$230 VGND VPWR sg13g2_decap_8
X$231 VGND VPWR sg13g2_decap_8
X$232 VGND VPWR sg13g2_decap_8
X$233 VGND VPWR sg13g2_decap_8
X$234 VGND VPWR sg13g2_decap_8
X$235 VGND VPWR sg13g2_decap_8
X$236 VGND VPWR sg13g2_decap_8
X$237 VGND VPWR sg13g2_decap_8
X$238 VGND VPWR sg13g2_decap_8
X$239 VGND VPWR sg13g2_decap_8
X$240 VGND VPWR sg13g2_decap_8
X$241 VGND VPWR sg13g2_decap_8
X$242 VGND VPWR sg13g2_decap_8
X$243 VGND VPWR sg13g2_decap_8
X$244 VGND VPWR sg13g2_decap_8
X$245 VGND VPWR sg13g2_decap_8
X$246 VGND VPWR sg13g2_decap_8
X$247 VGND VPWR sg13g2_decap_8
X$248 VGND VPWR sg13g2_decap_8
X$249 VGND VPWR sg13g2_decap_8
X$250 VGND VPWR sg13g2_decap_8
X$251 VGND VPWR sg13g2_decap_8
X$252 VGND VPWR sg13g2_decap_8
X$253 VGND VPWR sg13g2_decap_8
X$254 VGND VPWR sg13g2_decap_8
X$255 VGND VPWR sg13g2_decap_8
X$256 VGND VPWR sg13g2_decap_8
X$257 VGND VPWR sg13g2_decap_8
X$258 VGND VPWR sg13g2_decap_8
X$263 VGND VPWR sg13g2_decap_8
X$264 VGND VPWR sg13g2_decap_8
X$265 VGND VPWR sg13g2_decap_8
X$266 VGND VPWR sg13g2_decap_8
X$271 VGND VPWR sg13g2_decap_8
X$272 VGND VPWR sg13g2_decap_8
X$273 VGND VPWR sg13g2_decap_8
X$274 VGND VPWR sg13g2_decap_8
X$275 VGND VPWR sg13g2_decap_8
X$276 VGND VPWR sg13g2_decap_8
X$277 VGND VPWR sg13g2_decap_8
X$278 VGND VPWR sg13g2_decap_8
X$279 VGND VPWR sg13g2_decap_8
X$280 VGND VPWR sg13g2_decap_8
X$281 VGND VPWR sg13g2_decap_8
X$282 VGND VPWR sg13g2_decap_8
X$283 VGND VPWR sg13g2_decap_8
X$284 VGND VPWR sg13g2_decap_8
X$285 VGND VPWR sg13g2_decap_8
X$286 VGND VPWR sg13g2_decap_8
X$287 VGND VPWR sg13g2_decap_8
X$288 VGND VPWR sg13g2_decap_8
X$289 VGND VPWR sg13g2_decap_8
X$290 VGND VPWR sg13g2_decap_8
X$295 VGND VPWR sg13g2_decap_8
X$296 VGND VPWR sg13g2_decap_8
X$297 VGND VPWR sg13g2_decap_8
X$298 VGND VPWR sg13g2_decap_8
X$299 VGND VPWR sg13g2_decap_8
X$300 VGND VPWR sg13g2_decap_8
X$301 VGND VPWR sg13g2_decap_8
X$302 VGND VPWR sg13g2_decap_8
X$307 VGND VPWR sg13g2_decap_8
X$308 VGND VPWR sg13g2_decap_8
X$309 VGND VPWR sg13g2_decap_8
X$310 VGND VPWR sg13g2_decap_8
X$315 VGND VPWR sg13g2_decap_8
X$316 VGND VPWR sg13g2_decap_8
X$317 VGND VPWR sg13g2_decap_8
X$318 VGND VPWR sg13g2_decap_8
X$319 VGND VPWR sg13g2_decap_8
X$320 VGND VPWR sg13g2_decap_8
X$321 VGND VPWR sg13g2_decap_8
X$322 VGND VPWR sg13g2_decap_8
X$323 VGND VPWR sg13g2_decap_8
X$324 VGND VPWR sg13g2_decap_8
X$325 VGND VPWR sg13g2_decap_8
X$326 VGND VPWR sg13g2_decap_8
X$327 VGND VPWR sg13g2_decap_8
X$328 VGND VPWR sg13g2_decap_8
X$329 VGND VPWR sg13g2_decap_8
X$330 VGND VPWR sg13g2_decap_8
X$331 VGND VPWR sg13g2_decap_8
X$332 VGND VPWR sg13g2_decap_8
X$333 VGND VPWR sg13g2_decap_8
X$334 VGND VPWR sg13g2_decap_8
X$335 VGND VPWR sg13g2_decap_8
X$336 VGND VPWR sg13g2_decap_8
X$337 VGND VPWR sg13g2_decap_8
X$338 VGND VPWR sg13g2_decap_8
X$339 VGND VPWR sg13g2_decap_8
X$340 VGND VPWR sg13g2_decap_8
X$341 VGND VPWR sg13g2_decap_8
X$342 VGND VPWR sg13g2_decap_8
X$343 VGND VPWR sg13g2_decap_8
X$344 VGND VPWR sg13g2_decap_8
X$345 VGND VPWR sg13g2_decap_8
X$346 VGND VPWR sg13g2_decap_8
X$347 VGND VPWR sg13g2_decap_8
X$348 VGND VPWR sg13g2_decap_8
X$349 VGND VPWR sg13g2_decap_8
X$350 VGND VPWR sg13g2_decap_8
X$351 VGND VPWR sg13g2_decap_8
X$352 VGND VPWR sg13g2_decap_8
X$353 VGND VPWR sg13g2_decap_8
X$354 VGND VPWR sg13g2_decap_8
X$355 VGND VPWR sg13g2_decap_8
X$356 VGND VPWR sg13g2_decap_8
X$361 VGND VPWR sg13g2_decap_8
X$362 VGND VPWR sg13g2_decap_8
X$363 VGND VPWR sg13g2_decap_8
X$364 VGND VPWR sg13g2_decap_8
X$369 VGND VPWR sg13g2_decap_8
X$370 VGND VPWR sg13g2_decap_8
X$371 VGND VPWR sg13g2_decap_8
X$372 VGND VPWR sg13g2_decap_8
X$373 VGND VPWR sg13g2_decap_8
X$374 VGND VPWR sg13g2_decap_8
X$375 VGND VPWR sg13g2_decap_8
X$376 VGND VPWR sg13g2_decap_8
X$377 VGND VPWR sg13g2_decap_8
X$378 VGND VPWR sg13g2_decap_8
X$379 VGND VPWR sg13g2_decap_8
X$380 VGND VPWR sg13g2_decap_8
X$381 VGND VPWR sg13g2_decap_8
X$382 VGND VPWR sg13g2_decap_8
X$383 VGND VPWR sg13g2_decap_8
X$384 VGND VPWR sg13g2_decap_8
X$385 VGND VPWR sg13g2_decap_8
X$386 VGND VPWR sg13g2_decap_8
X$387 VGND VPWR sg13g2_decap_8
X$388 VGND VPWR sg13g2_decap_8
X$389 VGND VPWR sg13g2_decap_8
X$390 VGND VPWR sg13g2_decap_8
X$391 VGND VPWR sg13g2_decap_8
X$392 VGND VPWR sg13g2_decap_8
X$393 VGND VPWR sg13g2_decap_8
X$394 VGND VPWR sg13g2_decap_8
X$395 VGND VPWR sg13g2_decap_8
X$396 VGND VPWR sg13g2_decap_8
X$397 VGND VPWR sg13g2_decap_8
X$398 VGND VPWR sg13g2_decap_8
X$399 VGND VPWR sg13g2_decap_8
X$400 VGND VPWR sg13g2_decap_8
X$401 VGND VPWR sg13g2_decap_8
X$402 VGND VPWR sg13g2_decap_8
X$403 VGND VPWR sg13g2_decap_8
X$404 VGND VPWR sg13g2_decap_8
X$405 VGND VPWR sg13g2_decap_8
X$406 VGND VPWR sg13g2_decap_8
X$407 VGND VPWR sg13g2_decap_8
X$408 VGND VPWR sg13g2_decap_8
X$413 VGND VPWR sg13g2_decap_8
X$414 VGND VPWR sg13g2_decap_8
X$415 VGND VPWR sg13g2_decap_8
X$416 VGND VPWR sg13g2_decap_8
X$421 VGND VPWR sg13g2_decap_8
X$422 VGND VPWR sg13g2_decap_8
X$423 VGND VPWR sg13g2_decap_8
X$424 VGND VPWR sg13g2_decap_8
X$425 VGND VPWR sg13g2_decap_8
X$426 VGND VPWR sg13g2_decap_8
X$427 VGND VPWR sg13g2_decap_8
X$428 VGND VPWR sg13g2_decap_8
X$429 VGND VPWR sg13g2_decap_8
X$430 VGND VPWR sg13g2_decap_8
X$431 VGND VPWR sg13g2_decap_8
X$432 VGND VPWR sg13g2_decap_8
X$433 VGND VPWR sg13g2_decap_8
X$434 VGND VPWR sg13g2_decap_8
X$435 VGND VPWR sg13g2_decap_8
X$436 VGND VPWR sg13g2_decap_8
X$437 VGND VPWR sg13g2_decap_8
X$438 VGND VPWR sg13g2_decap_8
X$439 VGND VPWR sg13g2_decap_8
X$440 VGND VPWR sg13g2_decap_8
X$445 VGND VPWR sg13g2_decap_8
X$446 VGND VPWR sg13g2_decap_8
X$447 VGND VPWR sg13g2_decap_8
X$448 VGND VPWR sg13g2_decap_8
X$449 VGND VPWR sg13g2_decap_8
X$450 VGND VPWR sg13g2_decap_8
X$451 VGND VPWR sg13g2_decap_8
X$452 VGND VPWR sg13g2_decap_8
X$457 VGND VPWR sg13g2_decap_8
X$458 VGND VPWR sg13g2_decap_8
X$459 VGND VPWR sg13g2_decap_8
X$460 VGND VPWR sg13g2_decap_8
X$465 VGND VPWR sg13g2_decap_8
X$466 VGND VPWR sg13g2_decap_8
X$467 VGND VPWR sg13g2_decap_8
X$468 VGND VPWR sg13g2_decap_8
X$469 VGND VPWR sg13g2_decap_8
X$470 VGND VPWR sg13g2_decap_8
X$471 VGND VPWR sg13g2_decap_8
X$472 VGND VPWR sg13g2_decap_8
X$473 VGND VPWR sg13g2_decap_8
X$474 VGND VPWR sg13g2_decap_8
X$475 VGND VPWR sg13g2_decap_8
X$476 VGND VPWR sg13g2_decap_8
X$477 VGND VPWR sg13g2_decap_8
X$478 VGND VPWR sg13g2_decap_8
X$479 VGND VPWR sg13g2_decap_8
X$480 VGND VPWR sg13g2_decap_8
X$481 VGND VPWR sg13g2_decap_8
X$482 VGND VPWR sg13g2_decap_8
X$483 VGND VPWR sg13g2_decap_8
X$484 VGND VPWR sg13g2_decap_8
X$485 VGND VPWR sg13g2_decap_8
X$486 VGND VPWR sg13g2_decap_8
X$487 VGND VPWR sg13g2_decap_8
X$488 VGND VPWR sg13g2_decap_8
X$489 VGND VPWR sg13g2_decap_8
X$490 VGND VPWR sg13g2_decap_8
X$491 VGND VPWR sg13g2_decap_8
X$492 VGND VPWR sg13g2_decap_8
X$493 VGND VPWR sg13g2_decap_8
X$494 VGND VPWR sg13g2_decap_8
X$495 VGND VPWR sg13g2_decap_8
X$496 VGND VPWR sg13g2_decap_8
X$497 VGND VPWR sg13g2_decap_8
X$498 VGND VPWR sg13g2_decap_8
X$499 VGND VPWR sg13g2_decap_8
X$500 VGND VPWR sg13g2_decap_8
X$501 VGND VPWR sg13g2_decap_8
X$502 VGND VPWR sg13g2_decap_8
X$503 VGND VPWR sg13g2_decap_8
X$504 VGND VPWR sg13g2_decap_8
X$505 VGND VPWR sg13g2_decap_8
X$506 VGND VPWR sg13g2_decap_8
X$511 VGND VPWR sg13g2_decap_8
X$512 VGND VPWR sg13g2_decap_8
X$513 VGND VPWR sg13g2_decap_8
X$514 VGND VPWR sg13g2_decap_8
X$519 VGND VPWR sg13g2_decap_8
X$520 VGND VPWR sg13g2_decap_8
X$521 VGND VPWR sg13g2_decap_8
X$522 VGND VPWR sg13g2_decap_8
X$523 VGND VPWR sg13g2_decap_8
X$524 VGND VPWR sg13g2_decap_8
X$525 VGND VPWR sg13g2_decap_8
X$526 VGND VPWR sg13g2_decap_8
X$527 VGND VPWR sg13g2_decap_8
X$528 VGND VPWR sg13g2_decap_8
X$529 VGND VPWR sg13g2_decap_8
X$530 VGND VPWR sg13g2_decap_8
X$531 VGND VPWR sg13g2_decap_8
X$532 VGND VPWR sg13g2_decap_8
X$533 VGND VPWR sg13g2_decap_8
X$534 VGND VPWR sg13g2_decap_8
X$535 VGND VPWR sg13g2_decap_8
X$536 VGND VPWR sg13g2_decap_8
X$537 VGND VPWR sg13g2_decap_8
X$538 VGND VPWR sg13g2_decap_8
X$539 VGND VPWR sg13g2_decap_8
X$540 VGND VPWR sg13g2_decap_8
X$541 VGND VPWR sg13g2_decap_8
X$542 VGND VPWR sg13g2_decap_8
X$543 VGND VPWR sg13g2_decap_8
X$544 VGND VPWR sg13g2_decap_8
X$545 VGND VPWR sg13g2_decap_8
X$546 VGND VPWR sg13g2_decap_8
X$547 VGND VPWR sg13g2_decap_8
X$548 VGND VPWR sg13g2_decap_8
X$549 VGND VPWR sg13g2_decap_8
X$550 VGND VPWR sg13g2_decap_8
X$551 VGND VPWR sg13g2_decap_8
X$552 VGND VPWR sg13g2_decap_8
X$553 VGND VPWR sg13g2_decap_8
X$554 VGND VPWR sg13g2_decap_8
X$555 VGND VPWR sg13g2_decap_8
X$556 VGND VPWR sg13g2_decap_8
X$557 VGND VPWR sg13g2_decap_8
X$558 VGND VPWR sg13g2_decap_8
X$563 VGND VPWR sg13g2_decap_8
X$564 VGND VPWR sg13g2_decap_8
X$565 VGND VPWR sg13g2_decap_8
X$566 VGND VPWR sg13g2_decap_8
X$571 VGND VPWR sg13g2_decap_8
X$572 VGND VPWR sg13g2_decap_8
X$573 VGND VPWR sg13g2_decap_8
X$574 VGND VPWR sg13g2_decap_8
X$575 VGND VPWR sg13g2_decap_8
X$576 VGND VPWR sg13g2_decap_8
X$577 VGND VPWR sg13g2_decap_8
X$578 VGND VPWR sg13g2_decap_8
X$579 VGND VPWR sg13g2_decap_8
X$580 VGND VPWR sg13g2_decap_8
X$581 VGND VPWR sg13g2_decap_8
X$582 VGND VPWR sg13g2_decap_8
X$583 VGND VPWR sg13g2_decap_8
X$584 VGND VPWR sg13g2_decap_8
X$585 VGND VPWR sg13g2_decap_8
X$586 VGND VPWR sg13g2_decap_8
X$587 VGND VPWR sg13g2_decap_8
X$588 VGND VPWR sg13g2_decap_8
X$589 VGND VPWR sg13g2_decap_8
X$590 VGND VPWR sg13g2_decap_8
X$595 VGND VPWR sg13g2_decap_8
X$596 VGND VPWR sg13g2_decap_8
X$597 VGND VPWR sg13g2_decap_8
X$598 VGND VPWR sg13g2_decap_8
X$599 VGND VPWR sg13g2_decap_8
X$600 VGND VPWR sg13g2_decap_8
X$601 VGND VPWR sg13g2_decap_8
X$602 VGND VPWR sg13g2_decap_8
X$607 VGND VPWR sg13g2_decap_8
X$608 VGND VPWR sg13g2_decap_8
X$609 VGND VPWR sg13g2_decap_8
X$610 VGND VPWR sg13g2_decap_8
X$615 VGND VPWR sg13g2_decap_8
X$616 VGND VPWR sg13g2_decap_8
X$617 VGND VPWR sg13g2_decap_8
X$618 VGND VPWR sg13g2_decap_8
X$619 VGND VPWR sg13g2_decap_8
X$620 VGND VPWR sg13g2_decap_8
X$621 VGND VPWR sg13g2_decap_8
X$622 VGND VPWR sg13g2_decap_8
X$623 VGND VPWR sg13g2_decap_8
X$624 VGND VPWR sg13g2_decap_8
X$625 VGND VPWR sg13g2_decap_8
X$626 VGND VPWR sg13g2_decap_8
X$627 VGND VPWR sg13g2_decap_8
X$628 VGND VPWR sg13g2_decap_8
X$629 VGND VPWR sg13g2_decap_8
X$630 VGND VPWR sg13g2_decap_8
X$631 VGND VPWR sg13g2_decap_8
X$632 VGND VPWR sg13g2_decap_8
X$633 VGND VPWR sg13g2_decap_8
X$634 VGND VPWR sg13g2_decap_8
X$635 VGND VPWR sg13g2_decap_8
X$636 VGND VPWR sg13g2_decap_8
X$637 VGND VPWR sg13g2_decap_8
X$638 VGND VPWR sg13g2_decap_8
X$639 VGND VPWR sg13g2_decap_8
X$640 VGND VPWR sg13g2_decap_8
X$641 VGND VPWR sg13g2_decap_8
X$642 VGND VPWR sg13g2_decap_8
X$643 VGND VPWR sg13g2_decap_8
X$644 VGND VPWR sg13g2_decap_8
X$645 VGND VPWR sg13g2_decap_8
X$646 VGND VPWR sg13g2_decap_8
X$647 VGND VPWR sg13g2_decap_8
X$648 VGND VPWR sg13g2_decap_8
X$649 VGND VPWR sg13g2_decap_8
X$650 VGND VPWR sg13g2_decap_8
X$651 VGND VPWR sg13g2_decap_8
X$652 VGND VPWR sg13g2_decap_8
X$653 VGND VPWR sg13g2_decap_8
X$654 VGND VPWR sg13g2_decap_8
X$655 VGND VPWR sg13g2_decap_8
X$656 VGND VPWR sg13g2_decap_8
X$661 VGND VPWR sg13g2_decap_8
X$662 VGND VPWR sg13g2_decap_8
X$663 VGND VPWR sg13g2_decap_8
X$664 VGND VPWR sg13g2_decap_8
X$669 VGND VPWR sg13g2_decap_8
X$670 VGND VPWR sg13g2_decap_8
X$671 VGND VPWR sg13g2_decap_8
X$672 VGND VPWR sg13g2_decap_8
X$673 VGND VPWR sg13g2_decap_8
X$674 VGND VPWR sg13g2_decap_8
X$675 VGND VPWR sg13g2_decap_8
X$676 VGND VPWR sg13g2_decap_8
X$677 VGND VPWR sg13g2_decap_8
X$678 VGND VPWR sg13g2_decap_8
X$679 VGND VPWR sg13g2_decap_8
X$680 VGND VPWR sg13g2_decap_8
X$681 VGND VPWR sg13g2_decap_8
X$682 VGND VPWR sg13g2_decap_8
X$683 VGND VPWR sg13g2_decap_8
X$684 VGND VPWR sg13g2_decap_8
X$685 VGND VPWR sg13g2_decap_8
X$686 VGND VPWR sg13g2_decap_8
X$687 VGND VPWR sg13g2_decap_8
X$688 VGND VPWR sg13g2_decap_8
X$689 VGND VPWR sg13g2_decap_8
X$690 VGND VPWR sg13g2_decap_8
X$691 VGND VPWR sg13g2_decap_8
X$692 VGND VPWR sg13g2_decap_8
X$693 VGND VPWR sg13g2_decap_8
X$694 VGND VPWR sg13g2_decap_8
X$695 VGND VPWR sg13g2_decap_8
X$696 VGND VPWR sg13g2_decap_8
X$697 VGND VPWR sg13g2_decap_8
X$698 VGND VPWR sg13g2_decap_8
X$699 VGND VPWR sg13g2_decap_8
X$700 VGND VPWR sg13g2_decap_8
X$701 VGND VPWR sg13g2_decap_8
X$702 VGND VPWR sg13g2_decap_8
X$703 VGND VPWR sg13g2_decap_8
X$704 VGND VPWR sg13g2_decap_8
X$705 VGND VPWR sg13g2_decap_8
X$706 VGND VPWR sg13g2_decap_8
X$707 VGND VPWR sg13g2_decap_8
X$708 VGND VPWR sg13g2_decap_8
X$713 VGND VPWR sg13g2_decap_8
X$714 VGND VPWR sg13g2_decap_8
X$715 VGND VPWR sg13g2_decap_8
X$716 VGND VPWR sg13g2_decap_8
X$721 VGND VPWR sg13g2_decap_8
X$722 VGND VPWR sg13g2_decap_8
X$723 VGND VPWR sg13g2_decap_8
X$724 VGND VPWR sg13g2_decap_8
X$725 VGND VPWR sg13g2_decap_8
X$726 VGND VPWR sg13g2_decap_8
X$727 VGND VPWR sg13g2_decap_8
X$728 VGND VPWR sg13g2_decap_8
X$729 VGND VPWR sg13g2_decap_8
X$730 VGND VPWR sg13g2_decap_8
X$731 VGND VPWR sg13g2_decap_8
X$732 VGND VPWR sg13g2_decap_8
X$733 VGND VPWR sg13g2_decap_8
X$734 VGND VPWR sg13g2_decap_8
X$735 VGND VPWR sg13g2_decap_8
X$736 VGND VPWR sg13g2_decap_8
X$737 VGND VPWR sg13g2_decap_8
X$738 VGND VPWR sg13g2_decap_8
X$739 VGND VPWR sg13g2_decap_8
X$740 VGND VPWR sg13g2_decap_8
X$745 VGND VPWR sg13g2_decap_8
X$746 VGND VPWR sg13g2_decap_8
X$747 VGND VPWR sg13g2_decap_8
X$748 VGND VPWR sg13g2_decap_8
X$749 VGND VPWR sg13g2_decap_8
X$750 VGND VPWR sg13g2_decap_8
X$751 VGND VPWR sg13g2_decap_8
X$752 VGND VPWR sg13g2_decap_8
X$757 VGND VPWR sg13g2_decap_8
X$758 VGND VPWR sg13g2_decap_8
X$759 VGND VPWR sg13g2_decap_8
X$760 VGND VPWR sg13g2_decap_8
X$765 VGND VPWR sg13g2_decap_8
X$766 VGND VPWR sg13g2_decap_8
X$767 VGND VPWR sg13g2_decap_8
X$768 VGND VPWR sg13g2_decap_8
X$769 VGND VPWR sg13g2_decap_8
X$770 VGND VPWR sg13g2_decap_8
X$771 VGND VPWR sg13g2_decap_8
X$772 VGND VPWR sg13g2_decap_8
X$773 VGND VPWR sg13g2_decap_8
X$774 VGND VPWR sg13g2_decap_8
X$775 VGND VPWR sg13g2_decap_8
X$776 VGND VPWR sg13g2_decap_8
X$777 VGND VPWR sg13g2_decap_8
X$778 VGND VPWR sg13g2_decap_8
X$779 VGND VPWR sg13g2_decap_8
X$780 VGND VPWR sg13g2_decap_8
X$781 VGND VPWR sg13g2_decap_8
X$782 VGND VPWR sg13g2_decap_8
X$783 VGND VPWR sg13g2_decap_8
X$784 VGND VPWR sg13g2_decap_8
X$785 VGND VPWR sg13g2_decap_8
X$786 VGND VPWR sg13g2_decap_8
X$787 VGND VPWR sg13g2_decap_8
X$788 VGND VPWR sg13g2_decap_8
X$789 VGND VPWR sg13g2_decap_8
X$790 VGND VPWR sg13g2_decap_8
X$791 VGND VPWR sg13g2_decap_8
X$792 VGND VPWR sg13g2_decap_8
X$793 VGND VPWR sg13g2_decap_8
X$794 VGND VPWR sg13g2_decap_8
X$795 VGND VPWR sg13g2_decap_8
X$796 VGND VPWR sg13g2_decap_8
X$797 VGND VPWR sg13g2_decap_8
X$798 VGND VPWR sg13g2_decap_8
X$799 VGND VPWR sg13g2_decap_8
X$800 VGND VPWR sg13g2_decap_8
X$801 VGND VPWR sg13g2_decap_8
X$802 VGND VPWR sg13g2_decap_8
X$803 VGND VPWR sg13g2_decap_8
X$804 VGND VPWR sg13g2_decap_8
X$805 VGND VPWR sg13g2_decap_8
X$806 VGND VPWR sg13g2_decap_8
X$811 VGND VPWR sg13g2_decap_8
X$812 VGND VPWR sg13g2_decap_8
X$813 VGND VPWR sg13g2_decap_8
X$814 VGND VPWR sg13g2_decap_8
X$819 VGND VPWR sg13g2_decap_8
X$820 VGND VPWR sg13g2_decap_8
X$821 VGND VPWR sg13g2_decap_8
X$822 VGND VPWR sg13g2_decap_8
X$823 VGND VPWR sg13g2_decap_8
X$824 VGND VPWR sg13g2_decap_8
X$825 VGND VPWR sg13g2_decap_8
X$826 VGND VPWR sg13g2_decap_8
X$827 VGND VPWR sg13g2_decap_8
X$828 VGND VPWR sg13g2_decap_8
X$829 VGND VPWR sg13g2_decap_8
X$830 VGND VPWR sg13g2_decap_8
X$831 VGND VPWR sg13g2_decap_8
X$832 VGND VPWR sg13g2_decap_8
X$833 VGND VPWR sg13g2_decap_8
X$834 VGND VPWR sg13g2_decap_8
X$835 VGND VPWR sg13g2_decap_8
X$836 VGND VPWR sg13g2_decap_8
X$837 VGND VPWR sg13g2_decap_8
X$838 VGND VPWR sg13g2_decap_8
X$839 VGND VPWR sg13g2_decap_8
X$840 VGND VPWR sg13g2_decap_8
X$841 VGND VPWR sg13g2_decap_8
X$842 VGND VPWR sg13g2_decap_8
X$843 VGND VPWR sg13g2_decap_8
X$844 VGND VPWR sg13g2_decap_8
X$845 VGND VPWR sg13g2_decap_8
X$846 VGND VPWR sg13g2_decap_8
X$847 VGND VPWR sg13g2_decap_8
X$848 VGND VPWR sg13g2_decap_8
X$849 VGND VPWR sg13g2_decap_8
X$850 VGND VPWR sg13g2_decap_8
X$851 VGND VPWR sg13g2_decap_8
X$852 VGND VPWR sg13g2_decap_8
X$853 VGND VPWR sg13g2_decap_8
X$854 VGND VPWR sg13g2_decap_8
X$855 VGND VPWR sg13g2_decap_8
X$856 VGND VPWR sg13g2_decap_8
X$857 VGND VPWR sg13g2_decap_8
X$858 VGND VPWR sg13g2_decap_8
X$863 VGND VPWR sg13g2_decap_8
X$864 VGND VPWR sg13g2_decap_8
X$865 VGND VPWR sg13g2_decap_8
X$866 VGND VPWR sg13g2_decap_8
X$871 VGND VPWR sg13g2_decap_8
X$872 VGND VPWR sg13g2_decap_8
X$873 VGND VPWR sg13g2_decap_8
X$874 VGND VPWR sg13g2_decap_8
X$875 VGND VPWR sg13g2_decap_8
X$876 VGND VPWR sg13g2_decap_8
X$877 VGND VPWR sg13g2_decap_8
X$878 VGND VPWR sg13g2_decap_8
X$879 VGND VPWR sg13g2_decap_8
X$880 VGND VPWR sg13g2_decap_8
X$881 VGND VPWR sg13g2_decap_8
X$882 VGND VPWR sg13g2_decap_8
X$883 VGND VPWR sg13g2_decap_8
X$884 VGND VPWR sg13g2_decap_8
X$885 VGND VPWR sg13g2_decap_8
X$886 VGND VPWR sg13g2_decap_8
X$887 VGND VPWR sg13g2_decap_8
X$888 VGND VPWR sg13g2_decap_8
X$889 VGND VPWR sg13g2_decap_8
X$890 VGND VPWR sg13g2_decap_8
X$895 VGND VPWR sg13g2_decap_8
X$896 VGND VPWR sg13g2_decap_8
X$897 VGND VPWR sg13g2_decap_8
X$898 VGND VPWR sg13g2_decap_8
X$899 VGND VPWR sg13g2_decap_8
X$900 VGND VPWR sg13g2_decap_8
X$901 VGND VPWR sg13g2_decap_8
X$902 VGND VPWR sg13g2_decap_8
X$907 VGND VPWR sg13g2_decap_8
X$908 VGND VPWR sg13g2_decap_8
X$909 VGND VPWR sg13g2_decap_8
X$910 VGND VPWR sg13g2_decap_8
X$915 VGND VPWR sg13g2_decap_8
X$916 VGND VPWR sg13g2_decap_8
X$917 VGND VPWR sg13g2_decap_8
X$918 VGND VPWR sg13g2_decap_8
X$919 VGND VPWR sg13g2_decap_8
X$920 VGND VPWR sg13g2_decap_8
X$921 VGND VPWR sg13g2_decap_8
X$922 VGND VPWR sg13g2_decap_8
X$923 VGND VPWR sg13g2_decap_8
X$924 VGND VPWR sg13g2_decap_8
X$925 VGND VPWR sg13g2_decap_8
X$926 VGND VPWR sg13g2_decap_8
X$927 VGND VPWR sg13g2_decap_8
X$928 VGND VPWR sg13g2_decap_8
X$929 VGND VPWR sg13g2_decap_8
X$930 VGND VPWR sg13g2_decap_8
X$931 VGND VPWR sg13g2_decap_8
X$932 VGND VPWR sg13g2_decap_8
X$933 VGND VPWR sg13g2_decap_8
X$934 VGND VPWR sg13g2_decap_8
X$935 VGND VPWR sg13g2_decap_8
X$936 VGND VPWR sg13g2_decap_8
X$937 VGND VPWR sg13g2_decap_8
X$938 VGND VPWR sg13g2_decap_8
X$939 VGND VPWR sg13g2_decap_8
X$940 VGND VPWR sg13g2_decap_8
X$941 VGND VPWR sg13g2_decap_8
X$942 VGND VPWR sg13g2_decap_8
X$943 VGND VPWR sg13g2_decap_8
X$944 VGND VPWR sg13g2_decap_8
X$945 VGND VPWR sg13g2_decap_8
X$946 VGND VPWR sg13g2_decap_8
X$947 VGND VPWR sg13g2_decap_8
X$948 VGND VPWR sg13g2_decap_8
X$949 VGND VPWR sg13g2_decap_8
X$950 VGND VPWR sg13g2_decap_8
X$951 VGND VPWR sg13g2_decap_8
X$952 VGND VPWR sg13g2_decap_8
X$953 VGND VPWR sg13g2_decap_8
X$954 VGND VPWR sg13g2_decap_8
X$955 VGND VPWR sg13g2_decap_8
X$956 VGND VPWR sg13g2_decap_8
X$961 VGND VPWR sg13g2_decap_8
X$962 VGND VPWR sg13g2_decap_8
X$963 VGND VPWR sg13g2_decap_8
X$964 VGND VPWR sg13g2_decap_8
X$969 VGND VPWR sg13g2_decap_8
X$970 VGND VPWR sg13g2_decap_8
X$971 VGND VPWR sg13g2_decap_8
X$972 VGND VPWR sg13g2_decap_8
X$973 VGND VPWR sg13g2_decap_8
X$974 VGND VPWR sg13g2_decap_8
X$975 VGND VPWR sg13g2_decap_8
X$976 VGND VPWR sg13g2_decap_8
X$977 VGND VPWR sg13g2_decap_8
X$978 VGND VPWR sg13g2_decap_8
X$979 VGND VPWR sg13g2_decap_8
X$980 VGND VPWR sg13g2_decap_8
X$981 VGND VPWR sg13g2_decap_8
X$982 VGND VPWR sg13g2_decap_8
X$983 VGND VPWR sg13g2_decap_8
X$984 VGND VPWR sg13g2_decap_8
X$985 VGND VPWR sg13g2_decap_8
X$986 VGND VPWR sg13g2_decap_8
X$987 VGND VPWR sg13g2_decap_8
X$988 VGND VPWR sg13g2_decap_8
X$989 VGND VPWR sg13g2_decap_8
X$990 VGND VPWR sg13g2_decap_8
X$991 VGND VPWR sg13g2_decap_8
X$992 VGND VPWR sg13g2_decap_8
X$993 VGND VPWR sg13g2_decap_8
X$994 VGND VPWR sg13g2_decap_8
X$995 VGND VPWR sg13g2_decap_8
X$996 VGND VPWR sg13g2_decap_8
X$997 VGND VPWR sg13g2_decap_8
X$998 VGND VPWR sg13g2_decap_8
X$999 VGND VPWR sg13g2_decap_8
X$1000 VGND VPWR sg13g2_decap_8
X$1001 VGND VPWR sg13g2_decap_8
X$1002 VGND VPWR sg13g2_decap_8
X$1003 VGND VPWR sg13g2_decap_8
X$1004 VGND VPWR sg13g2_decap_8
X$1005 VGND VPWR sg13g2_decap_8
X$1006 VGND VPWR sg13g2_decap_8
X$1007 VGND VPWR sg13g2_decap_8
X$1008 VGND VPWR sg13g2_decap_8
X$1013 VGND VPWR sg13g2_decap_8
X$1014 VGND VPWR sg13g2_decap_8
X$1015 VGND VPWR sg13g2_decap_8
X$1016 VGND VPWR sg13g2_decap_8
X$1021 VGND VPWR sg13g2_decap_8
X$1022 VGND VPWR sg13g2_decap_8
X$1023 VGND VPWR sg13g2_decap_8
X$1024 VGND VPWR sg13g2_decap_8
X$1025 VGND VPWR sg13g2_decap_8
X$1026 VGND VPWR sg13g2_decap_8
X$1027 VGND VPWR sg13g2_decap_8
X$1028 VGND VPWR sg13g2_decap_8
X$1029 VGND VPWR sg13g2_decap_8
X$1030 VGND VPWR sg13g2_decap_8
X$1031 VGND VPWR sg13g2_decap_8
X$1032 VGND VPWR sg13g2_decap_8
X$1033 VGND VPWR sg13g2_decap_8
X$1034 VGND VPWR sg13g2_decap_8
X$1035 VGND VPWR sg13g2_decap_8
X$1036 VGND VPWR sg13g2_decap_8
X$1037 VGND VPWR sg13g2_decap_8
X$1038 VGND VPWR sg13g2_decap_8
X$1039 VGND VPWR sg13g2_decap_8
X$1040 VGND VPWR sg13g2_decap_8
X$1045 VGND VPWR sg13g2_decap_8
X$1046 VGND VPWR sg13g2_decap_8
X$1047 VGND VPWR sg13g2_decap_8
X$1048 VGND VPWR sg13g2_decap_8
X$1049 VGND VPWR sg13g2_decap_8
X$1050 VGND VPWR sg13g2_decap_8
X$1051 VGND VPWR sg13g2_decap_8
X$1052 VGND VPWR sg13g2_decap_8
X$1057 VGND VPWR sg13g2_decap_8
X$1058 VGND VPWR sg13g2_decap_8
X$1059 VGND VPWR sg13g2_decap_8
X$1060 VGND VPWR sg13g2_decap_8
X$1065 VGND VPWR sg13g2_decap_8
X$1066 VGND VPWR sg13g2_decap_8
X$1067 VGND VPWR sg13g2_decap_8
X$1068 VGND VPWR sg13g2_decap_8
X$1069 VGND VPWR sg13g2_decap_8
X$1070 VGND VPWR sg13g2_decap_8
X$1071 VGND VPWR sg13g2_decap_8
X$1072 VGND VPWR sg13g2_decap_8
X$1073 VGND VPWR sg13g2_decap_8
X$1074 VGND VPWR sg13g2_decap_8
X$1075 VGND VPWR sg13g2_decap_8
X$1076 VGND VPWR sg13g2_decap_8
X$1077 VGND VPWR sg13g2_decap_8
X$1078 VGND VPWR sg13g2_decap_8
X$1079 VGND VPWR sg13g2_decap_8
X$1080 VGND VPWR sg13g2_decap_8
X$1081 VGND VPWR sg13g2_decap_8
X$1082 VGND VPWR sg13g2_decap_8
X$1083 VGND VPWR sg13g2_decap_8
X$1084 VGND VPWR sg13g2_decap_8
X$1085 VGND VPWR sg13g2_decap_8
X$1086 VGND VPWR sg13g2_decap_8
X$1087 VGND VPWR sg13g2_decap_8
X$1088 VGND VPWR sg13g2_decap_8
X$1089 VGND VPWR sg13g2_decap_8
X$1090 VGND VPWR sg13g2_decap_8
X$1091 VGND VPWR sg13g2_decap_8
X$1092 VGND VPWR sg13g2_decap_8
X$1093 VGND VPWR sg13g2_decap_8
X$1094 VGND VPWR sg13g2_decap_8
X$1095 VGND VPWR sg13g2_decap_8
X$1096 VGND VPWR sg13g2_decap_8
X$1097 VGND VPWR sg13g2_decap_8
X$1098 VGND VPWR sg13g2_decap_8
X$1099 VGND VPWR sg13g2_decap_8
X$1100 VGND VPWR sg13g2_decap_8
X$1101 VGND VPWR sg13g2_decap_8
X$1102 VGND VPWR sg13g2_decap_8
X$1103 VGND VPWR sg13g2_decap_8
X$1104 VGND VPWR sg13g2_decap_8
X$1105 VGND VPWR sg13g2_decap_8
X$1106 VGND VPWR sg13g2_decap_8
X$1111 VGND VPWR sg13g2_decap_8
X$1112 VGND VPWR sg13g2_decap_8
X$1113 VGND VPWR sg13g2_decap_8
X$1114 VGND VPWR sg13g2_decap_8
X$1119 VGND VPWR sg13g2_decap_8
X$1120 VGND VPWR sg13g2_decap_8
X$1121 VGND VPWR sg13g2_decap_8
X$1122 VGND VPWR sg13g2_decap_8
X$1123 VGND VPWR sg13g2_decap_8
X$1124 VGND VPWR sg13g2_decap_8
X$1125 VGND VPWR sg13g2_decap_8
X$1126 VGND VPWR sg13g2_decap_8
X$1127 VGND VPWR sg13g2_decap_8
X$1128 VGND VPWR sg13g2_decap_8
X$1129 VGND VPWR sg13g2_decap_8
X$1130 VGND VPWR sg13g2_decap_8
X$1131 VGND VPWR sg13g2_decap_8
X$1132 VGND VPWR sg13g2_decap_8
X$1133 VGND VPWR sg13g2_decap_8
X$1134 VGND VPWR sg13g2_decap_8
X$1135 VGND VPWR sg13g2_decap_8
X$1136 VGND VPWR sg13g2_decap_8
X$1137 VGND VPWR sg13g2_decap_8
X$1138 VGND VPWR sg13g2_decap_8
X$1139 VGND VPWR sg13g2_decap_8
X$1140 VGND VPWR sg13g2_decap_8
X$1141 VGND VPWR sg13g2_decap_8
X$1142 VGND VPWR sg13g2_decap_8
X$1143 VGND VPWR sg13g2_decap_8
X$1144 VGND VPWR sg13g2_decap_8
X$1145 VGND VPWR sg13g2_decap_8
X$1146 VGND VPWR sg13g2_decap_8
X$1147 VGND VPWR sg13g2_decap_8
X$1148 VGND VPWR sg13g2_decap_8
X$1149 VGND VPWR sg13g2_decap_8
X$1150 VGND VPWR sg13g2_decap_8
X$1151 VGND VPWR sg13g2_decap_8
X$1152 VGND VPWR sg13g2_decap_8
X$1153 VGND VPWR sg13g2_decap_8
X$1154 VGND VPWR sg13g2_decap_8
X$1155 VGND VPWR sg13g2_decap_8
X$1156 VGND VPWR sg13g2_decap_8
X$1157 VGND VPWR sg13g2_decap_8
X$1158 VGND VPWR sg13g2_decap_8
X$1163 VGND VPWR sg13g2_decap_8
X$1164 VGND VPWR sg13g2_decap_8
X$1165 VGND VPWR sg13g2_decap_8
X$1166 VGND VPWR sg13g2_decap_8
X$1171 VGND VPWR sg13g2_decap_8
X$1172 VGND VPWR sg13g2_decap_8
X$1173 VGND VPWR sg13g2_decap_8
X$1174 VGND VPWR sg13g2_decap_8
X$1175 VGND VPWR sg13g2_decap_8
X$1176 VGND VPWR sg13g2_decap_8
X$1177 VGND VPWR sg13g2_decap_8
X$1178 VGND VPWR sg13g2_decap_8
X$1179 VGND VPWR sg13g2_decap_8
X$1180 VGND VPWR sg13g2_decap_8
X$1181 VGND VPWR sg13g2_decap_8
X$1182 VGND VPWR sg13g2_decap_8
X$1183 VGND VPWR sg13g2_decap_8
X$1184 VGND VPWR sg13g2_decap_8
X$1185 VGND VPWR sg13g2_decap_8
X$1186 VGND VPWR sg13g2_decap_8
X$1187 VGND VPWR sg13g2_decap_8
X$1188 VGND VPWR sg13g2_decap_8
X$1189 VGND VPWR sg13g2_decap_8
X$1190 VGND VPWR sg13g2_decap_8
X$1195 VGND VPWR sg13g2_decap_8
X$1196 VGND VPWR sg13g2_decap_8
X$1197 VGND VPWR sg13g2_decap_8
X$1198 VGND VPWR sg13g2_decap_8
X$1199 VGND VPWR sg13g2_decap_8
X$1200 VGND VPWR sg13g2_decap_8
X$1201 VGND VPWR sg13g2_decap_8
X$1202 VGND VPWR sg13g2_decap_8
X$1207 VGND VPWR sg13g2_decap_8
X$1208 VGND VPWR sg13g2_decap_8
X$1209 VGND VPWR sg13g2_decap_8
X$1210 VGND VPWR sg13g2_decap_8
X$1215 VGND VPWR sg13g2_decap_8
X$1216 VGND VPWR sg13g2_decap_8
X$1217 VGND VPWR sg13g2_decap_8
X$1218 VGND VPWR sg13g2_decap_8
X$1219 VGND VPWR sg13g2_decap_8
X$1220 VGND VPWR sg13g2_decap_8
X$1221 VGND VPWR sg13g2_decap_8
X$1222 VGND VPWR sg13g2_decap_8
X$1223 VGND VPWR sg13g2_decap_8
X$1224 VGND VPWR sg13g2_decap_8
X$1225 VGND VPWR sg13g2_decap_8
X$1226 VGND VPWR sg13g2_decap_8
X$1227 VGND VPWR sg13g2_decap_8
X$1228 VGND VPWR sg13g2_decap_8
X$1229 VGND VPWR sg13g2_decap_8
X$1230 VGND VPWR sg13g2_decap_8
X$1231 VGND VPWR sg13g2_decap_8
X$1232 VGND VPWR sg13g2_decap_8
X$1233 VGND VPWR sg13g2_decap_8
X$1234 VGND VPWR sg13g2_decap_8
X$1235 VGND VPWR sg13g2_decap_8
X$1236 VGND VPWR sg13g2_decap_8
X$1237 VGND VPWR sg13g2_decap_8
X$1238 VGND VPWR sg13g2_decap_8
X$1239 VGND VPWR sg13g2_decap_8
X$1240 VGND VPWR sg13g2_decap_8
X$1241 VGND VPWR sg13g2_decap_8
X$1242 VGND VPWR sg13g2_decap_8
X$1243 VGND VPWR sg13g2_decap_8
X$1244 VGND VPWR sg13g2_decap_8
X$1245 VGND VPWR sg13g2_decap_8
X$1246 VGND VPWR sg13g2_decap_8
X$1247 VGND VPWR sg13g2_decap_8
X$1248 VGND VPWR sg13g2_decap_8
X$1249 VGND VPWR sg13g2_decap_8
X$1250 VGND VPWR sg13g2_decap_8
X$1251 VGND VPWR sg13g2_decap_8
X$1252 VGND VPWR sg13g2_decap_8
X$1253 VGND VPWR sg13g2_decap_8
X$1254 VGND VPWR sg13g2_decap_8
X$1255 VGND VPWR sg13g2_decap_8
X$1256 VGND VPWR sg13g2_decap_8
X$1261 VGND VPWR sg13g2_decap_8
X$1262 VGND VPWR sg13g2_decap_8
X$1263 VGND VPWR sg13g2_decap_8
X$1264 VGND VPWR sg13g2_decap_8
X$1269 VGND VPWR sg13g2_decap_8
X$1270 VGND VPWR sg13g2_decap_8
X$1271 VGND VPWR sg13g2_decap_8
X$1272 VGND VPWR sg13g2_decap_8
X$1273 VGND VPWR sg13g2_decap_8
X$1274 VGND VPWR sg13g2_decap_8
X$1275 VGND VPWR sg13g2_decap_8
X$1276 VGND VPWR sg13g2_decap_8
X$1277 VGND VPWR sg13g2_decap_8
X$1278 VGND VPWR sg13g2_decap_8
X$1279 VGND VPWR sg13g2_decap_8
X$1280 VGND VPWR sg13g2_decap_8
X$1281 VGND VPWR sg13g2_decap_8
X$1282 VGND VPWR sg13g2_decap_8
X$1283 VGND VPWR sg13g2_decap_8
X$1284 VGND VPWR sg13g2_decap_8
X$1285 VGND VPWR sg13g2_decap_8
X$1286 VGND VPWR sg13g2_decap_8
X$1287 VGND VPWR sg13g2_decap_8
X$1288 VGND VPWR sg13g2_decap_8
X$1289 VGND VPWR sg13g2_decap_8
X$1290 VGND VPWR sg13g2_decap_8
X$1291 VGND VPWR sg13g2_decap_8
X$1292 VGND VPWR sg13g2_decap_8
X$1293 VGND VPWR sg13g2_decap_8
X$1294 VGND VPWR sg13g2_decap_8
X$1295 VGND VPWR sg13g2_decap_8
X$1296 VGND VPWR sg13g2_decap_8
X$1297 VGND VPWR sg13g2_decap_8
X$1298 VGND VPWR sg13g2_decap_8
X$1299 VGND VPWR sg13g2_decap_8
X$1300 VGND VPWR sg13g2_decap_8
X$1301 VGND VPWR sg13g2_decap_8
X$1302 VGND VPWR sg13g2_decap_8
X$1303 VGND VPWR sg13g2_decap_8
X$1304 VGND VPWR sg13g2_decap_8
X$1305 VGND VPWR sg13g2_decap_8
X$1306 VGND VPWR sg13g2_decap_8
X$1307 VGND VPWR sg13g2_decap_8
X$1308 VGND VPWR sg13g2_decap_8
X$1313 VGND VPWR sg13g2_decap_8
X$1314 VGND VPWR sg13g2_decap_8
X$1315 VGND VPWR sg13g2_decap_8
X$1316 VGND VPWR sg13g2_decap_8
X$1321 VGND VPWR sg13g2_decap_8
X$1322 VGND VPWR sg13g2_decap_8
X$1323 VGND VPWR sg13g2_decap_8
X$1324 VGND VPWR sg13g2_decap_8
X$1325 VGND VPWR sg13g2_decap_8
X$1326 VGND VPWR sg13g2_decap_8
X$1327 VGND VPWR sg13g2_decap_8
X$1328 VGND VPWR sg13g2_decap_8
X$1329 VGND VPWR sg13g2_decap_8
X$1330 VGND VPWR sg13g2_decap_8
X$1331 VGND VPWR sg13g2_decap_8
X$1332 VGND VPWR sg13g2_decap_8
X$1333 VGND VPWR sg13g2_decap_8
X$1334 VGND VPWR sg13g2_decap_8
X$1335 VGND VPWR sg13g2_decap_8
X$1336 VGND VPWR sg13g2_decap_8
X$1337 VGND VPWR sg13g2_decap_8
X$1338 VGND VPWR sg13g2_decap_8
X$1339 VGND VPWR sg13g2_decap_8
X$1340 VGND VPWR sg13g2_decap_8
X$1345 VGND VPWR sg13g2_decap_8
X$1346 VGND VPWR sg13g2_decap_8
X$1347 VGND VPWR sg13g2_decap_8
X$1348 VGND VPWR sg13g2_decap_8
X$1349 VGND VPWR sg13g2_decap_8
X$1350 VGND VPWR sg13g2_decap_8
X$1351 VGND VPWR sg13g2_decap_8
X$1352 VGND VPWR sg13g2_decap_8
X$1357 VGND VPWR sg13g2_decap_8
X$1358 VGND VPWR sg13g2_decap_8
X$1359 VGND VPWR sg13g2_decap_8
X$1360 VGND VPWR sg13g2_decap_8
X$1365 VGND VPWR sg13g2_decap_8
X$1366 VGND VPWR sg13g2_decap_8
X$1367 VGND VPWR sg13g2_decap_8
X$1368 VGND VPWR sg13g2_decap_8
X$1369 VGND VPWR sg13g2_decap_8
X$1370 VGND VPWR sg13g2_decap_8
X$1371 VGND VPWR sg13g2_decap_8
X$1372 VGND VPWR sg13g2_decap_8
X$1373 VGND VPWR sg13g2_decap_8
X$1374 VGND VPWR sg13g2_decap_8
X$1375 VGND VPWR sg13g2_decap_8
X$1376 VGND VPWR sg13g2_decap_8
X$1377 VGND VPWR sg13g2_decap_8
X$1378 VGND VPWR sg13g2_decap_8
X$1379 VGND VPWR sg13g2_decap_8
X$1380 VGND VPWR sg13g2_decap_8
X$1381 VGND VPWR sg13g2_decap_8
X$1382 VGND VPWR sg13g2_decap_8
X$1383 VGND VPWR sg13g2_decap_8
X$1384 VGND VPWR sg13g2_decap_8
X$1385 VGND VPWR sg13g2_decap_8
X$1386 VGND VPWR sg13g2_decap_8
X$1387 VGND VPWR sg13g2_decap_8
X$1388 VGND VPWR sg13g2_decap_8
X$1389 VGND VPWR sg13g2_decap_8
X$1390 VGND VPWR sg13g2_decap_8
X$1391 VGND VPWR sg13g2_decap_8
X$1392 VGND VPWR sg13g2_decap_8
X$1393 VGND VPWR sg13g2_decap_8
X$1394 VGND VPWR sg13g2_decap_8
X$1395 VGND VPWR sg13g2_decap_8
X$1396 VGND VPWR sg13g2_decap_8
X$1397 VGND VPWR sg13g2_decap_8
X$1398 VGND VPWR sg13g2_decap_8
X$1399 VGND VPWR sg13g2_decap_8
X$1400 VGND VPWR sg13g2_decap_8
X$1401 VGND VPWR sg13g2_decap_8
X$1402 VGND VPWR sg13g2_decap_8
X$1403 VGND VPWR sg13g2_decap_8
X$1404 VGND VPWR sg13g2_decap_8
X$1405 VGND VPWR sg13g2_decap_8
X$1406 VGND VPWR sg13g2_decap_8
X$1411 VGND VPWR sg13g2_decap_8
X$1412 VGND VPWR sg13g2_decap_8
X$1413 VGND VPWR sg13g2_decap_8
X$1414 VGND VPWR sg13g2_decap_8
X$1419 VGND VPWR sg13g2_decap_8
X$1420 VGND VPWR sg13g2_decap_8
X$1421 VGND VPWR sg13g2_decap_8
X$1422 VGND VPWR sg13g2_decap_8
X$1423 VGND VPWR sg13g2_decap_8
X$1424 VGND VPWR sg13g2_decap_8
X$1425 VGND VPWR sg13g2_decap_8
X$1426 VGND VPWR sg13g2_decap_8
X$1427 VGND VPWR sg13g2_decap_8
X$1428 VGND VPWR sg13g2_decap_8
X$1429 VGND VPWR sg13g2_decap_8
X$1430 VGND VPWR sg13g2_decap_8
X$1431 VGND VPWR sg13g2_decap_8
X$1432 VGND VPWR sg13g2_decap_8
X$1433 VGND VPWR sg13g2_decap_8
X$1434 VGND VPWR sg13g2_decap_8
X$1435 VGND VPWR sg13g2_decap_8
X$1436 VGND VPWR sg13g2_decap_8
X$1437 VGND VPWR sg13g2_decap_8
X$1438 VGND VPWR sg13g2_decap_8
X$1439 VGND VPWR sg13g2_decap_8
X$1440 VGND VPWR sg13g2_decap_8
X$1441 VGND VPWR sg13g2_decap_8
X$1442 VGND VPWR sg13g2_decap_8
X$1443 VGND VPWR sg13g2_decap_8
X$1444 VGND VPWR sg13g2_decap_8
X$1445 VGND VPWR sg13g2_decap_8
X$1446 VGND VPWR sg13g2_decap_8
X$1447 VGND VPWR sg13g2_decap_8
X$1448 VGND VPWR sg13g2_decap_8
X$1449 VGND VPWR sg13g2_decap_8
X$1450 VGND VPWR sg13g2_decap_8
X$1451 VGND VPWR sg13g2_decap_8
X$1452 VGND VPWR sg13g2_decap_8
X$1453 VGND VPWR sg13g2_decap_8
X$1454 VGND VPWR sg13g2_decap_8
X$1455 VGND VPWR sg13g2_decap_8
X$1456 VGND VPWR sg13g2_decap_8
X$1457 VGND VPWR sg13g2_decap_8
X$1458 VGND VPWR sg13g2_decap_8
X$1463 VGND VPWR sg13g2_decap_8
X$1464 VGND VPWR sg13g2_decap_8
X$1465 VGND VPWR sg13g2_decap_8
X$1466 VGND VPWR sg13g2_decap_8
X$1471 VGND VPWR sg13g2_decap_8
X$1472 VGND VPWR sg13g2_decap_8
X$1473 VGND VPWR sg13g2_decap_8
X$1474 VGND VPWR sg13g2_decap_8
X$1475 VGND VPWR sg13g2_decap_8
X$1476 VGND VPWR sg13g2_decap_8
X$1477 VGND VPWR sg13g2_decap_8
X$1478 VGND VPWR sg13g2_decap_8
X$1479 VGND VPWR sg13g2_decap_8
X$1480 VGND VPWR sg13g2_decap_8
X$1481 VGND VPWR sg13g2_decap_8
X$1482 VGND VPWR sg13g2_decap_8
X$1483 VGND VPWR sg13g2_decap_8
X$1484 VGND VPWR sg13g2_decap_8
X$1485 VGND VPWR sg13g2_decap_8
X$1486 VGND VPWR sg13g2_decap_8
X$1487 VGND VPWR sg13g2_decap_8
X$1488 VGND VPWR sg13g2_decap_8
X$1489 VGND VPWR sg13g2_decap_8
X$1490 VGND VPWR sg13g2_decap_8
X$1495 VGND VPWR sg13g2_decap_8
X$1496 VGND VPWR sg13g2_decap_8
X$1497 VGND VPWR sg13g2_decap_8
X$1498 VGND VPWR sg13g2_decap_8
X$1499 VGND VPWR sg13g2_decap_8
X$1500 VGND VPWR sg13g2_decap_8
X$1501 VGND VPWR sg13g2_decap_8
X$1502 VGND VPWR sg13g2_decap_8
X$1507 VGND VPWR sg13g2_decap_8
X$1508 VGND VPWR sg13g2_decap_8
X$1509 VGND VPWR sg13g2_decap_8
X$1510 VGND VPWR sg13g2_decap_8
X$1515 VGND VPWR sg13g2_decap_8
X$1516 VGND VPWR sg13g2_decap_8
X$1517 VGND VPWR sg13g2_decap_8
X$1518 VGND VPWR sg13g2_decap_8
X$1519 VGND VPWR sg13g2_decap_8
X$1520 VGND VPWR sg13g2_decap_8
X$1521 VGND VPWR sg13g2_decap_8
X$1522 VGND VPWR sg13g2_decap_8
X$1523 VGND VPWR sg13g2_decap_8
X$1524 VGND VPWR sg13g2_decap_8
X$1525 VGND VPWR sg13g2_decap_8
X$1526 VGND VPWR sg13g2_decap_8
X$1527 VGND VPWR sg13g2_decap_8
X$1528 VGND VPWR sg13g2_decap_8
X$1529 VGND VPWR sg13g2_decap_8
X$1530 VGND VPWR sg13g2_decap_8
X$1531 VGND VPWR sg13g2_decap_8
X$1532 VGND VPWR sg13g2_decap_8
X$1533 VGND VPWR sg13g2_decap_8
X$1534 VGND VPWR sg13g2_decap_8
X$1535 VGND VPWR sg13g2_decap_8
X$1536 VGND VPWR sg13g2_decap_8
X$1537 VGND VPWR sg13g2_decap_8
X$1538 VGND VPWR sg13g2_decap_8
X$1539 VGND VPWR sg13g2_decap_8
X$1540 VGND VPWR sg13g2_decap_8
X$1541 VGND VPWR sg13g2_decap_8
X$1542 VGND VPWR sg13g2_decap_8
X$1543 VGND VPWR sg13g2_decap_8
X$1544 VGND VPWR sg13g2_decap_8
X$1545 VGND VPWR sg13g2_decap_8
X$1546 VGND VPWR sg13g2_decap_8
X$1547 VGND VPWR sg13g2_decap_8
X$1548 VGND VPWR sg13g2_decap_8
X$1549 VGND VPWR sg13g2_decap_8
X$1550 VGND VPWR sg13g2_decap_8
X$1551 VGND VPWR sg13g2_decap_8
X$1552 VGND VPWR sg13g2_decap_8
X$1553 VGND VPWR sg13g2_decap_8
X$1554 VGND VPWR sg13g2_decap_8
X$1555 VGND VPWR sg13g2_decap_8
X$1556 VGND VPWR sg13g2_decap_8
X$1561 VGND VPWR sg13g2_decap_8
X$1562 VGND VPWR sg13g2_decap_8
X$1563 VGND VPWR sg13g2_decap_8
X$1564 VGND VPWR sg13g2_decap_8
X$1569 VGND VPWR sg13g2_decap_8
X$1570 VGND VPWR sg13g2_decap_8
X$1571 VGND VPWR sg13g2_decap_8
X$1572 VGND VPWR sg13g2_decap_8
X$1573 VGND VPWR sg13g2_decap_8
X$1574 VGND VPWR sg13g2_decap_8
X$1575 VGND VPWR sg13g2_decap_8
X$1576 VGND VPWR sg13g2_decap_8
X$1577 VGND VPWR sg13g2_decap_8
X$1578 VGND VPWR sg13g2_decap_8
X$1579 VGND VPWR sg13g2_decap_8
X$1580 VGND VPWR sg13g2_decap_8
X$1581 VGND VPWR sg13g2_decap_8
X$1582 VGND VPWR sg13g2_decap_8
X$1583 VGND VPWR sg13g2_decap_8
X$1584 VGND VPWR sg13g2_decap_8
X$1585 VGND VPWR sg13g2_decap_8
X$1586 VGND VPWR sg13g2_decap_8
X$1587 VGND VPWR sg13g2_decap_8
X$1588 VGND VPWR sg13g2_decap_8
X$1589 VGND VPWR sg13g2_decap_8
X$1590 VGND VPWR sg13g2_decap_8
X$1591 VGND VPWR sg13g2_decap_8
X$1592 VGND VPWR sg13g2_decap_8
X$1593 VGND VPWR sg13g2_decap_8
X$1594 VGND VPWR sg13g2_decap_8
X$1595 VGND VPWR sg13g2_decap_8
X$1596 VGND VPWR sg13g2_decap_8
X$1597 VGND VPWR sg13g2_decap_8
X$1598 VGND VPWR sg13g2_decap_8
X$1599 VGND VPWR sg13g2_decap_8
X$1600 VGND VPWR sg13g2_decap_8
X$1601 VGND VPWR sg13g2_decap_8
X$1602 VGND VPWR sg13g2_decap_8
X$1603 VGND VPWR sg13g2_decap_8
X$1604 VGND VPWR sg13g2_decap_8
X$1605 VGND VPWR sg13g2_decap_8
X$1606 VGND VPWR sg13g2_decap_8
X$1607 VGND VPWR sg13g2_decap_8
X$1608 VGND VPWR sg13g2_decap_8
X$1613 VGND VPWR sg13g2_decap_8
X$1614 VGND VPWR sg13g2_decap_8
X$1615 VGND VPWR sg13g2_decap_8
X$1616 VGND VPWR sg13g2_decap_8
X$1621 VGND VPWR sg13g2_decap_8
X$1622 VGND VPWR sg13g2_decap_8
X$1623 VGND VPWR sg13g2_decap_8
X$1624 VGND VPWR sg13g2_decap_8
X$1625 VGND VPWR sg13g2_decap_8
X$1626 VGND VPWR sg13g2_decap_8
X$1627 VGND VPWR sg13g2_decap_8
X$1628 VGND VPWR sg13g2_decap_8
X$1629 VGND VPWR sg13g2_decap_8
X$1630 VGND VPWR sg13g2_decap_8
X$1631 VGND VPWR sg13g2_decap_8
X$1632 VGND VPWR sg13g2_decap_8
X$1633 VGND VPWR sg13g2_decap_8
X$1634 VGND VPWR sg13g2_decap_8
X$1635 VGND VPWR sg13g2_decap_8
X$1636 VGND VPWR sg13g2_decap_8
X$1637 VGND VPWR sg13g2_decap_8
X$1638 VGND VPWR sg13g2_decap_8
X$1639 VGND VPWR sg13g2_decap_8
X$1640 VGND VPWR sg13g2_decap_8
X$1645 VGND VPWR sg13g2_decap_8
X$1646 VGND VPWR sg13g2_decap_8
X$1647 VGND VPWR sg13g2_decap_8
X$1648 VGND VPWR sg13g2_decap_8
X$1649 VGND VPWR sg13g2_decap_8
X$1650 VGND VPWR sg13g2_decap_8
X$1651 VGND VPWR sg13g2_decap_8
X$1652 VGND VPWR sg13g2_decap_8
X$1657 VGND VPWR sg13g2_decap_8
X$1658 VGND VPWR sg13g2_decap_8
X$1659 VGND VPWR sg13g2_decap_8
X$1660 VGND VPWR sg13g2_decap_8
X$1665 VGND VPWR sg13g2_decap_8
X$1666 VGND VPWR sg13g2_decap_8
X$1667 VGND VPWR sg13g2_decap_8
X$1668 VGND VPWR sg13g2_decap_8
X$1669 VGND VPWR sg13g2_decap_8
X$1670 VGND VPWR sg13g2_decap_8
X$1671 VGND VPWR sg13g2_decap_8
X$1672 VGND VPWR sg13g2_decap_8
X$1673 VGND VPWR sg13g2_decap_8
X$1674 VGND VPWR sg13g2_decap_8
X$1675 VGND VPWR sg13g2_decap_8
X$1676 VGND VPWR sg13g2_decap_8
X$1677 VGND VPWR sg13g2_decap_8
X$1678 VGND VPWR sg13g2_decap_8
X$1679 VGND VPWR sg13g2_decap_8
X$1680 VGND VPWR sg13g2_decap_8
X$1681 VGND VPWR sg13g2_decap_8
X$1682 VGND VPWR sg13g2_decap_8
X$1683 VGND VPWR sg13g2_decap_8
X$1684 VGND VPWR sg13g2_decap_8
X$1685 VGND VPWR sg13g2_decap_8
X$1686 VGND VPWR sg13g2_decap_8
X$1687 VGND VPWR sg13g2_decap_8
X$1688 VGND VPWR sg13g2_decap_8
X$1689 VGND VPWR sg13g2_decap_8
X$1690 VGND VPWR sg13g2_decap_8
X$1691 VGND VPWR sg13g2_decap_8
X$1692 VGND VPWR sg13g2_decap_8
X$1693 VGND VPWR sg13g2_decap_8
X$1694 VGND VPWR sg13g2_decap_8
X$1695 VGND VPWR sg13g2_decap_8
X$1696 VGND VPWR sg13g2_decap_8
X$1697 VGND VPWR sg13g2_decap_8
X$1698 VGND VPWR sg13g2_decap_8
X$1699 VGND VPWR sg13g2_decap_8
X$1700 VGND VPWR sg13g2_decap_8
X$1701 VGND VPWR sg13g2_decap_8
X$1702 VGND VPWR sg13g2_decap_8
X$1703 VGND VPWR sg13g2_decap_8
X$1704 VGND VPWR sg13g2_decap_8
X$1705 VGND VPWR sg13g2_decap_8
X$1706 VGND VPWR sg13g2_decap_8
X$1711 VGND VPWR sg13g2_decap_8
X$1712 VGND VPWR sg13g2_decap_8
X$1713 VGND VPWR sg13g2_decap_8
X$1714 VGND VPWR sg13g2_decap_8
X$1719 VGND VPWR sg13g2_decap_8
X$1720 VGND VPWR sg13g2_decap_8
X$1721 VGND VPWR sg13g2_decap_8
X$1722 VGND VPWR sg13g2_decap_8
X$1723 VGND VPWR sg13g2_decap_8
X$1724 VGND VPWR sg13g2_decap_8
X$1725 VGND VPWR sg13g2_decap_8
X$1726 VGND VPWR sg13g2_decap_8
X$1727 VGND VPWR sg13g2_decap_8
X$1728 VGND VPWR sg13g2_decap_8
X$1729 VGND VPWR sg13g2_decap_8
X$1730 VGND VPWR sg13g2_decap_8
X$1731 VGND VPWR sg13g2_decap_8
X$1732 VGND VPWR sg13g2_decap_8
X$1733 VGND VPWR sg13g2_decap_8
X$1734 VGND VPWR sg13g2_decap_8
X$1735 VGND VPWR sg13g2_decap_8
X$1736 VGND VPWR sg13g2_decap_8
X$1737 VGND VPWR sg13g2_decap_8
X$1738 VGND VPWR sg13g2_decap_8
X$1739 VGND VPWR sg13g2_decap_8
X$1740 VGND VPWR sg13g2_decap_8
X$1741 VGND VPWR sg13g2_decap_8
X$1742 VGND VPWR sg13g2_decap_8
X$1743 VGND VPWR sg13g2_decap_8
X$1744 VGND VPWR sg13g2_decap_8
X$1745 VGND VPWR sg13g2_decap_8
X$1746 VGND VPWR sg13g2_decap_8
X$1747 VGND VPWR sg13g2_decap_8
X$1748 VGND VPWR sg13g2_decap_8
X$1749 VGND VPWR sg13g2_decap_8
X$1750 VGND VPWR sg13g2_decap_8
X$1751 VGND VPWR sg13g2_decap_8
X$1752 VGND VPWR sg13g2_decap_8
X$1753 VGND VPWR sg13g2_decap_8
X$1754 VGND VPWR sg13g2_decap_8
X$1755 VGND VPWR sg13g2_decap_8
X$1756 VGND VPWR sg13g2_decap_8
X$1757 VGND VPWR sg13g2_decap_8
X$1758 VGND VPWR sg13g2_decap_8
X$1763 VGND VPWR sg13g2_decap_8
X$1764 VGND VPWR sg13g2_decap_8
X$1765 VGND VPWR sg13g2_decap_8
X$1766 VGND VPWR sg13g2_decap_8
X$1771 VGND VPWR sg13g2_decap_8
X$1772 VGND VPWR sg13g2_decap_8
X$1773 VGND VPWR sg13g2_decap_8
X$1774 VGND VPWR sg13g2_decap_8
X$1775 VGND VPWR sg13g2_decap_8
X$1776 VGND VPWR sg13g2_decap_8
X$1777 VGND VPWR sg13g2_decap_8
X$1778 VGND VPWR sg13g2_decap_8
X$1779 VGND VPWR sg13g2_decap_8
X$1780 VGND VPWR sg13g2_decap_8
X$1781 VGND VPWR sg13g2_decap_8
X$1782 VGND VPWR sg13g2_decap_8
X$1783 VGND VPWR sg13g2_decap_8
X$1784 VGND VPWR sg13g2_decap_8
X$1785 VGND VPWR sg13g2_decap_8
X$1786 VGND VPWR sg13g2_decap_8
X$1787 VGND VPWR sg13g2_decap_8
X$1788 VGND VPWR sg13g2_decap_8
X$1789 VGND VPWR sg13g2_decap_8
X$1790 VGND VPWR sg13g2_decap_8
X$1795 VGND VPWR sg13g2_decap_8
X$1796 VGND VPWR sg13g2_decap_8
X$1797 VGND VPWR sg13g2_decap_8
X$1798 VGND VPWR sg13g2_decap_8
X$1799 VGND VPWR sg13g2_decap_8
X$1800 VGND VPWR sg13g2_decap_8
X$1801 VGND VPWR sg13g2_decap_8
X$1802 VGND VPWR sg13g2_decap_8
X$1807 VGND VPWR sg13g2_decap_8
X$1808 VGND VPWR sg13g2_decap_8
X$1809 VGND VPWR sg13g2_decap_8
X$1810 VGND VPWR sg13g2_decap_8
X$1815 VGND VPWR sg13g2_decap_8
X$1816 VGND VPWR sg13g2_decap_8
X$1817 VGND VPWR sg13g2_decap_8
X$1818 VGND VPWR sg13g2_decap_8
X$1819 VGND VPWR sg13g2_decap_8
X$1820 VGND VPWR sg13g2_decap_8
X$1821 VGND VPWR sg13g2_decap_8
X$1822 VGND VPWR sg13g2_decap_8
X$1823 VGND VPWR sg13g2_decap_8
X$1824 VGND VPWR sg13g2_decap_8
X$1825 VGND VPWR sg13g2_decap_8
X$1826 VGND VPWR sg13g2_decap_8
X$1827 VGND VPWR sg13g2_decap_8
X$1828 VGND VPWR sg13g2_decap_8
X$1829 VGND VPWR sg13g2_decap_8
X$1830 VGND VPWR sg13g2_decap_8
X$1831 VGND VPWR sg13g2_decap_8
X$1832 VGND VPWR sg13g2_decap_8
X$1833 VGND VPWR sg13g2_decap_8
X$1834 VGND VPWR sg13g2_decap_8
X$1835 VGND VPWR sg13g2_decap_8
X$1836 VGND VPWR sg13g2_decap_8
X$1837 VGND VPWR sg13g2_decap_8
X$1838 VGND VPWR sg13g2_decap_8
X$1839 VGND VPWR sg13g2_decap_8
X$1840 VGND VPWR sg13g2_decap_8
X$1841 VGND VPWR sg13g2_decap_8
X$1842 VGND VPWR sg13g2_decap_8
X$1843 VGND VPWR sg13g2_decap_8
X$1844 VGND VPWR sg13g2_decap_8
X$1845 VGND VPWR sg13g2_decap_8
X$1846 VGND VPWR sg13g2_decap_8
X$1847 VGND VPWR sg13g2_decap_8
X$1848 VGND VPWR sg13g2_decap_8
X$1849 VGND VPWR sg13g2_decap_8
X$1850 VGND VPWR sg13g2_decap_8
X$1851 VGND VPWR sg13g2_decap_8
X$1852 VGND VPWR sg13g2_decap_8
X$1853 VGND VPWR sg13g2_decap_8
X$1854 VGND VPWR sg13g2_decap_8
X$1855 VGND VPWR sg13g2_decap_8
X$1856 VGND VPWR sg13g2_decap_8
X$1861 VGND VPWR sg13g2_decap_8
X$1862 VGND VPWR sg13g2_decap_8
X$1863 VGND VPWR sg13g2_decap_8
X$1864 VGND VPWR sg13g2_decap_8
X$1869 VGND VPWR sg13g2_decap_8
X$1870 VGND VPWR sg13g2_decap_8
X$1871 VGND VPWR sg13g2_decap_8
X$1872 VGND VPWR sg13g2_decap_8
X$1873 VGND VPWR sg13g2_decap_8
X$1874 VGND VPWR sg13g2_decap_8
X$1875 VGND VPWR sg13g2_decap_8
X$1876 VGND VPWR sg13g2_decap_8
X$1877 VGND VPWR sg13g2_decap_8
X$1878 VGND VPWR sg13g2_decap_8
X$1879 VGND VPWR sg13g2_decap_8
X$1880 VGND VPWR sg13g2_decap_8
X$1881 VGND VPWR sg13g2_decap_8
X$1882 VGND VPWR sg13g2_decap_8
X$1883 VGND VPWR sg13g2_decap_8
X$1884 VGND VPWR sg13g2_decap_8
X$1885 VGND VPWR sg13g2_decap_8
X$1886 VGND VPWR sg13g2_decap_8
X$1887 VGND VPWR sg13g2_decap_8
X$1888 VGND VPWR sg13g2_decap_8
X$1889 VGND VPWR sg13g2_decap_8
X$1890 VGND VPWR sg13g2_decap_8
X$1891 VGND VPWR sg13g2_decap_8
X$1892 VGND VPWR sg13g2_decap_8
X$1893 VGND VPWR sg13g2_decap_8
X$1894 VGND VPWR sg13g2_decap_8
X$1895 VGND VPWR sg13g2_decap_8
X$1896 VGND VPWR sg13g2_decap_8
X$1897 VGND VPWR sg13g2_decap_8
X$1898 VGND VPWR sg13g2_decap_8
X$1899 VGND VPWR sg13g2_decap_8
X$1900 VGND VPWR sg13g2_decap_8
X$1901 VGND VPWR sg13g2_decap_8
X$1902 VGND VPWR sg13g2_decap_8
X$1903 VGND VPWR sg13g2_decap_8
X$1904 VGND VPWR sg13g2_decap_8
X$1905 VGND VPWR sg13g2_decap_8
X$1906 VGND VPWR sg13g2_decap_8
X$1907 VGND VPWR sg13g2_decap_8
X$1908 VGND VPWR sg13g2_decap_8
X$1913 VGND VPWR sg13g2_decap_8
X$1914 VGND VPWR sg13g2_decap_8
X$1915 VGND VPWR sg13g2_decap_8
X$1916 VGND VPWR sg13g2_decap_8
X$1921 VGND VPWR sg13g2_decap_8
X$1922 VGND VPWR sg13g2_decap_8
X$1923 VGND VPWR sg13g2_decap_8
X$1924 VGND VPWR sg13g2_decap_8
X$1925 VGND VPWR sg13g2_decap_8
X$1926 VGND VPWR sg13g2_decap_8
X$1927 VGND VPWR sg13g2_decap_8
X$1928 VGND VPWR sg13g2_decap_8
X$1929 VGND VPWR sg13g2_decap_8
X$1930 VGND VPWR sg13g2_decap_8
X$1931 VGND VPWR sg13g2_decap_8
X$1932 VGND VPWR sg13g2_decap_8
X$1933 VGND VPWR sg13g2_decap_8
X$1934 VGND VPWR sg13g2_decap_8
X$1935 VGND VPWR sg13g2_decap_8
X$1936 VGND VPWR sg13g2_decap_8
X$1937 VGND VPWR sg13g2_decap_8
X$1938 VGND VPWR sg13g2_decap_8
X$1939 VGND VPWR sg13g2_decap_8
X$1940 VGND VPWR sg13g2_decap_8
X$1945 VGND VPWR sg13g2_decap_8
X$1946 VGND VPWR sg13g2_decap_8
X$1947 VGND VPWR sg13g2_decap_8
X$1948 VGND VPWR sg13g2_decap_8
X$1949 VGND VPWR sg13g2_decap_8
X$1950 VGND VPWR sg13g2_decap_8
X$1951 VGND VPWR sg13g2_decap_8
X$1952 VGND VPWR sg13g2_decap_8
X$1957 VGND VPWR sg13g2_decap_8
X$1958 VGND VPWR sg13g2_decap_8
X$1959 VGND VPWR sg13g2_decap_8
X$1960 VGND VPWR sg13g2_decap_8
X$1965 VGND VPWR sg13g2_decap_8
X$1966 VGND VPWR sg13g2_decap_8
X$1967 VGND VPWR sg13g2_decap_8
X$1968 VGND VPWR sg13g2_decap_8
X$1969 VGND VPWR sg13g2_decap_8
X$1970 VGND VPWR sg13g2_decap_8
X$1971 VGND VPWR sg13g2_decap_8
X$1972 VGND VPWR sg13g2_decap_8
X$1973 VGND VPWR sg13g2_decap_8
X$1974 VGND VPWR sg13g2_decap_8
X$1975 VGND VPWR sg13g2_decap_8
X$1976 VGND VPWR sg13g2_decap_8
X$1977 VGND VPWR sg13g2_decap_8
X$1978 VGND VPWR sg13g2_decap_8
X$1979 VGND VPWR sg13g2_decap_8
X$1980 VGND VPWR sg13g2_decap_8
X$1981 VGND VPWR sg13g2_decap_8
X$1982 VGND VPWR sg13g2_decap_8
X$1983 VGND VPWR sg13g2_decap_8
X$1984 VGND VPWR sg13g2_decap_8
X$1985 VGND VPWR sg13g2_decap_8
X$1986 VGND VPWR sg13g2_decap_8
X$1987 VGND VPWR sg13g2_decap_8
X$1988 VGND VPWR sg13g2_decap_8
X$1989 VGND VPWR sg13g2_decap_8
X$1990 VGND VPWR sg13g2_decap_8
X$1991 VGND VPWR sg13g2_decap_8
X$1992 VGND VPWR sg13g2_decap_8
X$1993 VGND VPWR sg13g2_decap_8
X$1994 VGND VPWR sg13g2_decap_8
X$1995 VGND VPWR sg13g2_decap_8
X$1996 VGND VPWR sg13g2_decap_8
X$1997 VGND VPWR sg13g2_decap_8
X$1998 VGND VPWR sg13g2_decap_8
X$1999 VGND VPWR sg13g2_decap_8
X$2000 VGND VPWR sg13g2_decap_8
X$2001 VGND VPWR sg13g2_decap_8
X$2002 VGND VPWR sg13g2_decap_8
X$2003 VGND VPWR sg13g2_decap_8
X$2004 VGND VPWR sg13g2_decap_8
X$2005 VGND VPWR sg13g2_decap_8
X$2006 VGND VPWR sg13g2_decap_8
X$2011 VGND VPWR sg13g2_decap_8
X$2012 VGND VPWR sg13g2_decap_8
X$2013 VGND VPWR sg13g2_decap_8
X$2014 VGND VPWR sg13g2_decap_8
X$2019 VGND VPWR sg13g2_decap_8
X$2020 VGND VPWR sg13g2_decap_8
X$2021 VGND VPWR sg13g2_decap_8
X$2022 VGND VPWR sg13g2_decap_8
X$2023 VGND VPWR sg13g2_decap_8
X$2024 VGND VPWR sg13g2_decap_8
X$2025 VGND VPWR sg13g2_decap_8
X$2026 VGND VPWR sg13g2_decap_8
X$2027 VGND VPWR sg13g2_decap_8
X$2028 VGND VPWR sg13g2_decap_8
X$2029 VGND VPWR sg13g2_decap_8
X$2030 VGND VPWR sg13g2_decap_8
X$2031 VGND VPWR sg13g2_decap_8
X$2032 VGND VPWR sg13g2_decap_8
X$2033 VGND VPWR sg13g2_decap_8
X$2034 VGND VPWR sg13g2_decap_8
X$2035 VGND VPWR sg13g2_decap_8
X$2036 VGND VPWR sg13g2_decap_8
X$2037 VGND VPWR sg13g2_decap_8
X$2038 VGND VPWR sg13g2_decap_8
X$2039 VGND VPWR sg13g2_decap_8
X$2040 VGND VPWR sg13g2_decap_8
X$2041 VGND VPWR sg13g2_decap_8
X$2042 VGND VPWR sg13g2_decap_8
X$2043 VGND VPWR sg13g2_decap_8
X$2044 VGND VPWR sg13g2_decap_8
X$2045 VGND VPWR sg13g2_decap_8
X$2046 VGND VPWR sg13g2_decap_8
X$2047 VGND VPWR sg13g2_decap_8
X$2048 VGND VPWR sg13g2_decap_8
X$2049 VGND VPWR sg13g2_decap_8
X$2050 VGND VPWR sg13g2_decap_8
X$2051 VGND VPWR sg13g2_decap_8
X$2052 VGND VPWR sg13g2_decap_8
X$2053 VGND VPWR sg13g2_decap_8
X$2054 VGND VPWR sg13g2_decap_8
X$2055 VGND VPWR sg13g2_decap_8
X$2056 VGND VPWR sg13g2_decap_8
X$2057 VGND VPWR sg13g2_decap_8
X$2058 VGND VPWR sg13g2_decap_8
X$2063 VGND VPWR sg13g2_decap_8
X$2064 VGND VPWR sg13g2_decap_8
X$2065 VGND VPWR sg13g2_decap_8
X$2066 VGND VPWR sg13g2_decap_8
X$2071 VGND VPWR sg13g2_decap_8
X$2072 VGND VPWR sg13g2_decap_8
X$2073 VGND VPWR sg13g2_decap_8
X$2074 VGND VPWR sg13g2_decap_8
X$2075 VGND VPWR sg13g2_decap_8
X$2076 VGND VPWR sg13g2_decap_8
X$2077 VGND VPWR sg13g2_decap_8
X$2078 VGND VPWR sg13g2_decap_8
X$2079 VGND VPWR sg13g2_decap_8
X$2080 VGND VPWR sg13g2_decap_8
X$2081 VGND VPWR sg13g2_decap_8
X$2082 VGND VPWR sg13g2_decap_8
X$2083 VGND VPWR sg13g2_decap_8
X$2084 VGND VPWR sg13g2_decap_8
X$2085 VGND VPWR sg13g2_decap_8
X$2086 VGND VPWR sg13g2_decap_8
X$2087 VGND VPWR sg13g2_decap_8
X$2088 VGND VPWR sg13g2_decap_8
X$2089 VGND VPWR sg13g2_decap_8
X$2090 VGND VPWR sg13g2_decap_8
X$2095 VGND VPWR sg13g2_decap_8
X$2096 VGND VPWR sg13g2_decap_8
X$2097 VGND VPWR sg13g2_decap_8
X$2098 VGND VPWR sg13g2_decap_8
X$2099 VGND VPWR sg13g2_decap_8
X$2100 VGND VPWR sg13g2_decap_8
X$2101 VGND VPWR sg13g2_decap_8
X$2102 VGND VPWR sg13g2_decap_8
X$2107 VGND VPWR sg13g2_decap_8
X$2108 VGND VPWR sg13g2_decap_8
X$2109 VGND VPWR sg13g2_decap_8
X$2110 VGND VPWR sg13g2_decap_8
X$2115 VGND VPWR sg13g2_decap_8
X$2116 VGND VPWR sg13g2_decap_8
X$2117 VGND VPWR sg13g2_decap_8
X$2118 VGND VPWR sg13g2_decap_8
X$2119 VGND VPWR sg13g2_decap_8
X$2120 VGND VPWR sg13g2_decap_8
X$2121 VGND VPWR sg13g2_decap_8
X$2122 VGND VPWR sg13g2_decap_8
X$2123 VGND VPWR sg13g2_decap_8
X$2124 VGND VPWR sg13g2_decap_8
X$2125 VGND VPWR sg13g2_decap_8
X$2126 VGND VPWR sg13g2_decap_8
X$2127 VGND VPWR sg13g2_decap_8
X$2128 VGND VPWR sg13g2_decap_8
X$2129 VGND VPWR sg13g2_decap_8
X$2130 VGND VPWR sg13g2_decap_8
X$2131 VGND VPWR sg13g2_decap_8
X$2132 VGND VPWR sg13g2_decap_8
X$2133 VGND VPWR sg13g2_decap_8
X$2134 VGND VPWR sg13g2_decap_8
X$2135 VGND VPWR sg13g2_decap_8
X$2136 VGND VPWR sg13g2_decap_8
X$2137 VGND VPWR sg13g2_decap_8
X$2138 VGND VPWR sg13g2_decap_8
X$2139 VGND VPWR sg13g2_decap_8
X$2140 VGND VPWR sg13g2_decap_8
X$2141 VGND VPWR sg13g2_decap_8
X$2142 VGND VPWR sg13g2_decap_8
X$2143 VGND VPWR sg13g2_decap_8
X$2144 VGND VPWR sg13g2_decap_8
X$2145 VGND VPWR sg13g2_decap_8
X$2146 VGND VPWR sg13g2_decap_8
X$2147 VGND VPWR sg13g2_decap_8
X$2148 VGND VPWR sg13g2_decap_8
X$2149 VGND VPWR sg13g2_decap_8
X$2150 VGND VPWR sg13g2_decap_8
X$2151 VGND VPWR sg13g2_decap_8
X$2152 VGND VPWR sg13g2_decap_8
X$2153 VGND VPWR sg13g2_decap_8
X$2154 VGND VPWR sg13g2_decap_8
X$2155 VGND VPWR sg13g2_decap_8
X$2156 VGND VPWR sg13g2_decap_8
X$2161 VGND VPWR sg13g2_decap_8
X$2162 VGND VPWR sg13g2_decap_8
X$2163 VGND VPWR sg13g2_decap_8
X$2164 VGND VPWR sg13g2_decap_8
X$2169 VGND VPWR sg13g2_decap_8
X$2170 VGND VPWR sg13g2_decap_8
X$2171 VGND VPWR sg13g2_decap_8
X$2172 VGND VPWR sg13g2_decap_8
X$2173 VGND VPWR sg13g2_decap_8
X$2174 VGND VPWR sg13g2_decap_8
X$2175 VGND VPWR sg13g2_decap_8
X$2176 VGND VPWR sg13g2_decap_8
X$2177 VGND VPWR sg13g2_decap_8
X$2178 VGND VPWR sg13g2_decap_8
X$2179 VGND VPWR sg13g2_decap_8
X$2180 VGND VPWR sg13g2_decap_8
X$2181 VGND VPWR sg13g2_decap_8
X$2183 VGND ui_in[4] \$35 ui_in[3] \$44 VPWR sg13g2_a21oi_1
X$2184 VGND \$46 \$51 \$35 VPWR sg13g2_nand2_1
X$2185 VGND VPWR sg13g2_decap_8
X$2186 VGND VPWR sg13g2_decap_8
X$2187 VGND VPWR sg13g2_decap_8
X$2189 VGND \$49 \$57 ui_in[0] VPWR sg13g2_nand2_1
X$2190 VGND VPWR sg13g2_decap_8
X$2191 VGND VPWR sg13g2_decap_8
X$2192 VGND VPWR sg13g2_decap_8
X$2193 VGND VPWR sg13g2_decap_8
X$2194 VGND VPWR sg13g2_decap_8
X$2195 VGND VPWR sg13g2_decap_8
X$2196 VGND VPWR sg13g2_decap_8
X$2197 VGND VPWR sg13g2_decap_8
X$2198 VGND VPWR sg13g2_decap_8
X$2199 VGND VPWR sg13g2_decap_8
X$2200 VGND VPWR sg13g2_decap_8
X$2201 VGND VPWR sg13g2_decap_8
X$2202 VGND VPWR sg13g2_decap_8
X$2203 VGND VPWR sg13g2_decap_8
X$2204 VGND VPWR sg13g2_decap_8
X$2205 VGND VPWR sg13g2_decap_8
X$2206 VGND VPWR sg13g2_decap_8
X$2207 VGND VPWR sg13g2_decap_4
X$2209 VGND VPWR sg13g2_decap_8
X$2210 VGND ui_in[3] \$56 \$38 VPWR sg13g2_nor2_1
X$2211 VGND VPWR sg13g2_decap_8
X$2212 VGND VPWR sg13g2_decap_8
X$2213 VGND VPWR sg13g2_decap_8
X$2218 VGND VPWR sg13g2_decap_8
X$2219 VGND VPWR sg13g2_decap_8
X$2220 VGND VPWR sg13g2_decap_8
X$2221 VGND VPWR sg13g2_decap_8
X$2226 VGND VPWR sg13g2_decap_8
X$2227 VGND VPWR sg13g2_decap_8
X$2228 VGND VPWR sg13g2_decap_8
X$2229 VGND VPWR sg13g2_decap_8
X$2230 VGND VPWR sg13g2_decap_8
X$2231 VGND VPWR sg13g2_decap_8
X$2232 VGND VPWR sg13g2_decap_8
X$2233 VGND VPWR sg13g2_decap_8
X$2234 VGND VPWR sg13g2_decap_8
X$2235 VGND VPWR sg13g2_decap_8
X$2236 VGND VPWR sg13g2_decap_8
X$2237 VGND VPWR sg13g2_decap_8
X$2238 VGND VPWR sg13g2_decap_8
X$2239 VGND VPWR sg13g2_decap_8
X$2240 VGND VPWR sg13g2_decap_8
X$2241 VGND VPWR sg13g2_decap_8
X$2242 VGND VPWR sg13g2_decap_8
X$2243 VGND VPWR sg13g2_decap_8
X$2244 VGND VPWR sg13g2_decap_8
X$2245 VGND VPWR sg13g2_decap_4
X$2249 VGND VPWR sg13g2_decap_8
X$2250 VGND VPWR sg13g2_decap_8
X$2251 VGND VPWR sg13g2_decap_8
X$2252 VGND VPWR sg13g2_decap_8
X$2257 VGND VPWR sg13g2_decap_8
X$2258 VGND VPWR sg13g2_decap_8
X$2263 VGND VPWR sg13g2_decap_8
X$2264 VGND VPWR sg13g2_decap_8
X$2265 VGND VPWR sg13g2_decap_8
X$2266 VGND VPWR sg13g2_decap_8
X$2267 VGND VPWR sg13g2_decap_8
X$2268 VGND VPWR sg13g2_decap_8
X$2269 VGND VPWR sg13g2_decap_8
X$2270 VGND VPWR sg13g2_decap_8
X$2271 VGND VPWR sg13g2_decap_8
X$2272 VGND VPWR sg13g2_decap_8
X$2273 VGND VPWR sg13g2_decap_8
X$2274 VGND VPWR sg13g2_decap_8
X$2275 VGND VPWR sg13g2_decap_8
X$2276 VGND VPWR sg13g2_decap_8
X$2277 VGND VPWR sg13g2_decap_8
X$2278 VGND VPWR sg13g2_decap_8
X$2279 VGND VPWR sg13g2_decap_8
X$2280 VGND VPWR sg13g2_decap_8
X$2281 VGND VPWR sg13g2_decap_8
X$2282 VGND VPWR sg13g2_decap_8
X$2283 VGND VPWR sg13g2_decap_8
X$2288 VGND VPWR sg13g2_decap_8
X$2289 VGND VPWR sg13g2_decap_8
X$2294 VGND VPWR sg13g2_decap_8
X$2296 VGND ui_in[1] ui_in[0] \$58 VPWR sg13g2_xor2_1
X$2300 VGND ui_in[2] \$58 \$68 VPWR sg13g2_xor2_1
X$2303 VGND \$56 \$60 \$68 VPWR sg13g2_and2_1
X$2305 VGND \$151 \$56 \$68 ui_in[4] VPWR sg13g2_o21ai_1
X$2307 VGND \$111 \$60 \$151 \$51 VPWR sg13g2_o21ai_1
X$2310 VGND ui_in[3] \$58 \$46 \$49 VPWR sg13g2_nand3b_1
X$2320 VGND ui_in[1] \$44 ui_in[2] VPWR sg13g2_nor2b_1
X$2328 VGND ui_in[2] \$49 ui_in[1] VPWR sg13g2_nand2b_1
X$2332 VGND \$162 ui_in[3] \$57 \$35 VPWR sg13g2_o21ai_1
X$2336 VGND ui_in[3] \$63 \$57 VPWR sg13g2_nand2b_1
X$2339 VGND VPWR sg13g2_decap_8
X$2341 VGND VPWR sg13g2_decap_4
X$2342 VGND \$178 \$72 \$56 \$52 VPWR sg13g2_nor3_1
X$2343 VGND ui_in[1] \$72 \$92 VPWR sg13g2_nor2_1
X$2345 VGND VPWR sg13g2_decap_4
X$2347 VGND \$125 ui_in[1] ui_in[0] ui_in[3] VPWR sg13g2_o21ai_1
X$2349 VGND ui_in[0] \$92 ui_in[2] VPWR sg13g2_or2_1
X$2351 VGND ui_in[3] \$64 ui_in[1] VPWR sg13g2_nand2b_1
X$2354 VGND ui_in[2] \$52 ui_in[1] VPWR sg13g2_and2_1
X$2358 VGND ui_in[0] \$65 ui_in[3] VPWR sg13g2_nand2b_1
X$2361 VGND \$64 \$65 ui_in[2] \$131 VPWR sg13g2_nand3_1
X$2370 VGND \$56 \$79 \$98 VPWR sg13g2_nand2b_1
X$2374 VGND ui_in[4] \$98 ui_in[3] \$38 VPWR sg13g2_a21oi_1
X$2381 VGND \$67 \$131 ui_in[4] \$148 VPWR sg13g2_nand3_1
X$2382 VGND ui_in[2] \$38 ui_in[1] VPWR sg13g2_nor2_1
X$2385 VGND VPWR sg13g2_decap_4
X$2391 VGND ui_in[1] \$78 ui_in[0] VPWR sg13g2_nor2b_1
X$2392 VGND \$78 \$67 ui_in[3] \$100 VPWR sg13g2_a21oi_1
X$2395 VGND VPWR sg13g2_decap_8
X$2396 VGND VPWR sg13g2_decap_8
X$2397 VGND VPWR sg13g2_decap_8
X$2398 VGND VPWR sg13g2_decap_8
X$2399 VGND VPWR sg13g2_decap_8
X$2400 VGND VPWR sg13g2_decap_8
X$2401 VGND VPWR sg13g2_decap_8
X$2402 VGND VPWR sg13g2_decap_8
X$2403 VGND VPWR sg13g2_decap_4
X$2514 VGND VPWR sg13g2_decap_8
X$2515 VGND VPWR sg13g2_decap_8
X$2516 VGND VPWR sg13g2_decap_8
X$2517 VGND VPWR sg13g2_decap_8
X$2519 VGND VPWR sg13g2_decap_8
X$2520 VGND VPWR sg13g2_decap_8
X$2521 VGND VPWR sg13g2_decap_8
X$2522 VGND VPWR sg13g2_decap_8
X$2523 VGND VPWR sg13g2_decap_8
X$2524 VGND VPWR sg13g2_decap_8
X$2525 VGND VPWR sg13g2_decap_8
X$2526 VGND VPWR sg13g2_decap_8
X$2527 VGND VPWR sg13g2_decap_8
X$2528 VGND VPWR sg13g2_decap_8
X$2529 VGND VPWR sg13g2_decap_8
X$2530 VGND VPWR sg13g2_decap_8
X$2531 VGND VPWR sg13g2_decap_8
X$2532 VGND VPWR sg13g2_decap_8
X$2533 VGND VPWR sg13g2_decap_8
X$2534 VGND VPWR sg13g2_decap_8
X$2535 VGND VPWR sg13g2_decap_8
X$2536 VGND VPWR sg13g2_decap_8
X$2537 VGND VPWR sg13g2_decap_8
X$2538 VGND VPWR sg13g2_decap_8
X$2539 VGND VPWR sg13g2_decap_8
X$2540 VGND VPWR sg13g2_decap_8
X$2541 VGND VPWR sg13g2_decap_8
X$2543 VGND VPWR sg13g2_decap_8
X$2544 VGND VPWR sg13g2_decap_8
X$2545 VGND VPWR sg13g2_decap_4
X$2546 VGND ui_in[0] \$197 ui_in[1] VPWR sg13g2_nand2b_1
X$2547 VGND ui_in[3] \$105 ui_in[2] ui_in[1] VPWR sg13g2_a21oi_1
X$2548 VGND VPWR sg13g2_decap_4
X$2549 VGND \$200 ui_in[2] \$58 \$105 VPWR sg13g2_o21ai_1
X$2550 VGND VPWR sg13g2_decap_4
X$2552 VGND ui_in[4] \$110 ui_in[5] VPWR sg13g2_nor2b_1
X$2555 VGND VPWR sg13g2_decap_8
X$2559 VGND \$58 \$92 \$105 \$157 VPWR sg13g2_a21o_1
X$2562 VGND VPWR sg13g2_decap_8
X$2564 VGND VPWR sg13g2_decap_8
X$2565 VGND \$162 \$181 ui_in[5] \$208 VPWR sg13g2_nand3_1
X$2566 VGND \$185 \$63 \$110 \$182 VPWR sg13g2_nand3_1
X$2569 VGND \$105 \$124 \$92 VPWR sg13g2_nand2_1
X$2570 VGND \$125 \$38 \$100 \$185 VPWR sg13g2_or3_1
X$2572 VGND \$187 \$135 \$125 \$124 VPWR sg13g2_o21ai_1
X$2573 VGND VPWR sg13g2_decap_8
X$2577 VGND \$189 \$100 \$125 ui_in[4] VPWR sg13g2_o21ai_1
X$2581 VGND VPWR sg13g2_decap_8
X$2585 VGND VPWR sg13g2_decap_8
X$2586 VGND VPWR sg13g2_decap_8
X$2588 VGND VPWR sg13g2_decap_4
X$2590 VGND \$148 \$79 ui_in[5] \$222 VPWR sg13g2_nand3_1
X$2592 VGND VPWR sg13g2_decap_8
X$2595 VGND VPWR sg13g2_decap_4
X$2597 VGND \$133 \$192 \$181 ui_in[4] VPWR sg13g2_nand3b_1
X$2598 VGND \$133 \$135 \$78 ui_in[3] VPWR sg13g2_nor3_1
X$2600 VGND ui_in[2] \$100 ui_in[0] VPWR sg13g2_nor2_1
X$2602 VGND VPWR sg13g2_decap_8
X$2603 VGND VPWR sg13g2_decap_8
X$2604 VGND VPWR sg13g2_decap_8
X$2605 VGND VPWR sg13g2_decap_8
X$2606 VGND VPWR sg13g2_decap_8
X$2607 VGND VPWR sg13g2_decap_8
X$2608 VGND VPWR sg13g2_decap_8
X$2609 VGND VPWR sg13g2_decap_8
X$2612 VGND VPWR sg13g2_decap_8
X$2613 VGND VPWR sg13g2_decap_8
X$2614 VGND VPWR sg13g2_decap_8
X$2615 VGND VPWR sg13g2_decap_8
X$2619 VGND VPWR sg13g2_decap_8
X$2620 VGND VPWR sg13g2_decap_8
X$2622 VGND VPWR sg13g2_decap_8
X$2623 VGND VPWR sg13g2_decap_8
X$2624 VGND VPWR sg13g2_decap_8
X$2625 VGND VPWR sg13g2_decap_8
X$2626 VGND VPWR sg13g2_decap_8
X$2627 VGND VPWR sg13g2_decap_8
X$2628 VGND VPWR sg13g2_decap_8
X$2629 VGND VPWR sg13g2_decap_8
X$2630 VGND VPWR sg13g2_decap_8
X$2631 VGND VPWR sg13g2_decap_8
X$2632 VGND VPWR sg13g2_decap_8
X$2633 VGND VPWR sg13g2_decap_8
X$2634 VGND VPWR sg13g2_decap_8
X$2635 VGND VPWR sg13g2_decap_8
X$2636 VGND VPWR sg13g2_decap_8
X$2637 VGND VPWR sg13g2_decap_8
X$2638 VGND VPWR sg13g2_decap_8
X$2639 VGND VPWR sg13g2_decap_8
X$2640 VGND VPWR sg13g2_decap_8
X$2641 VGND VPWR sg13g2_decap_8
X$2642 VGND VPWR sg13g2_decap_8
X$2646 VGND VPWR sg13g2_decap_8
X$2647 VGND VPWR sg13g2_decap_8
X$2649 VGND VPWR sg13g2_decap_4
X$2651 VGND \$100 \$305 ui_in[2] \$58 VPWR sg13g2_a21oi_1
X$2657 VGND \$197 ui_in[2] ui_in[3] \$257 VPWR sg13g2_nand3_1
X$2668 VGND VPWR sg13g2_decap_4
X$2671 VGND \$257 \$200 \$110 \$354 VPWR sg13g2_nand3_1
X$2679 VGND VPWR sg13g2_decap_8
X$2683 VGND VPWR sg13g2_decap_8
X$2686 VGND VPWR sg13g2_decap_4
X$2689 VGND \$291 \$58 ui_in[2] \$365 VPWR sg13g2_or3_1
X$2698 VGND \$264 ui_in[3] \$306 \$157 VPWR sg13g2_o21ai_1
X$2700 VGND ui_in[6] \$265 \$249 \$264 VPWR sg13g2_a21oi_1
X$2702 VGND \$227 ui_in[7] \$228 \$182 \$208 \$265 VPWR sg13g2_a221oi_1
X$2712 VGND VPWR sg13g2_decap_8
X$2722 VGND VPWR sg13g2_decap_8
X$2732 VGND \$228 \$296 \$248 \$268 \$249 \$187 VPWR sg13g2_a221oi_1
X$2745 VGND \$229 \$271 \$178 \$249 VPWR sg13g2_o21ai_1
X$2748 VGND VPWR sg13g2_decap_4
X$2750 VGND \$64 \$323 \$92 \$253 VPWR sg13g2_a21oi_1
X$2760 VGND \$253 \$274 \$92 \$329 VPWR sg13g2_nand3_1
X$2762 VGND ui_in[4] \$232 \$52 VPWR sg13g2_nor2b_1
X$2764 VGND \$335 ui_in[5] \$232 \$334 \$276 \$329 VPWR sg13g2_a221oi_1
X$2766 VGND \$65 \$334 ui_in[2] VPWR sg13g2_nand2_1
X$2768 VGND VPWR sg13g2_decap_8
X$2774 VGND VPWR sg13g2_decap_8
X$2782 VGND VPWR sg13g2_decap_8
X$2784 VGND VPWR sg13g2_decap_4
X$2789 VGND ui_in[0] \$135 ui_in[2] VPWR sg13g2_nor2b_1
X$2796 VGND \$283 \$253 ui_in[3] \$192 VPWR sg13g2_nand3_1
X$2807 VGND ui_in[0] \$253 ui_in[2] VPWR sg13g2_nand2_1
X$2811 VGND VPWR sg13g2_decap_8
X$2812 VGND VPWR sg13g2_decap_8
X$2813 VGND VPWR sg13g2_decap_8
X$2814 VGND VPWR sg13g2_decap_8
X$2815 VGND VPWR sg13g2_decap_8
X$2816 VGND VPWR sg13g2_decap_8
X$2817 VGND VPWR sg13g2_decap_8
X$2818 VGND VPWR sg13g2_decap_8
X$2978 VGND VPWR sg13g2_decap_8
X$2979 VGND VPWR sg13g2_decap_8
X$2980 VGND VPWR sg13g2_decap_8
X$2981 VGND VPWR sg13g2_decap_8
X$2986 VGND VPWR sg13g2_decap_8
X$2987 VGND VPWR sg13g2_decap_8
X$2988 VGND VPWR sg13g2_decap_8
X$2989 VGND VPWR sg13g2_decap_8
X$2990 VGND VPWR sg13g2_decap_8
X$2991 VGND VPWR sg13g2_decap_8
X$2992 VGND VPWR sg13g2_decap_8
X$2993 VGND VPWR sg13g2_decap_8
X$2994 VGND VPWR sg13g2_decap_8
X$2995 VGND VPWR sg13g2_decap_8
X$2996 VGND VPWR sg13g2_decap_8
X$2997 VGND VPWR sg13g2_decap_8
X$2998 VGND VPWR sg13g2_decap_8
X$2999 VGND VPWR sg13g2_decap_8
X$3000 VGND VPWR sg13g2_decap_8
X$3001 VGND VPWR sg13g2_decap_8
X$3002 VGND VPWR sg13g2_decap_8
X$3003 VGND VPWR sg13g2_decap_8
X$3004 VGND VPWR sg13g2_decap_8
X$3005 VGND VPWR sg13g2_decap_8
X$3006 VGND VPWR sg13g2_decap_8
X$3007 VGND VPWR sg13g2_decap_8
X$3008 VGND VPWR sg13g2_decap_8
X$3013 VGND VPWR sg13g2_decap_8
X$3014 VGND VPWR sg13g2_decap_8
X$3015 VGND \$197 \$310 ui_in[3] VPWR sg13g2_nand2_1
X$3016 VGND \$105 \$311 \$306 VPWR sg13g2_nand2_1
X$3017 VGND \$197 \$253 \$306 ui_in[3] VPWR \$414 sg13g2_nand4_1
X$3018 VGND \$357 \$38 \$310 \$311 VPWR sg13g2_o21ai_1
X$3019 VGND VPWR sg13g2_decap_8
X$3020 VGND VPWR sg13g2_decap_8
X$3021 VGND VPWR sg13g2_decap_4
X$3023 VGND ui_in[3] \$291 \$248 VPWR sg13g2_nand2b_1
X$3024 VGND \$419 \$291 \$315 ui_in[6] VPWR sg13g2_o21ai_1
X$3026 VGND \$135 \$315 \$44 VPWR sg13g2_nor2_1
X$3027 VGND VPWR sg13g2_decap_8
X$3028 VGND VPWR sg13g2_decap_4
X$3030 VGND \$365 \$318 \$229 ui_in[6] VPWR \$382 sg13g2_nand4_1
X$3031 VGND \$63 \$384 \$110 \$318 VPWR sg13g2_nand3_1
X$3032 VGND VPWR sg13g2_decap_4
X$3033 VGND \$248 \$105 \$306 \$386 VPWR sg13g2_nand3_1
X$3035 VGND VPWR sg13g2_decap_4
X$3037 VGND \$274 \$268 \$411 VPWR sg13g2_and2_1
X$3038 VGND VPWR sg13g2_decap_8
X$3039 VGND VPWR sg13g2_decap_8
X$3040 VGND VPWR sg13g2_decap_8
X$3042 VGND \$336 \$283 \$291 \$100 VPWR sg13g2_nor3_1
X$3044 VGND \$410 \$335 \$336 \$296 VPWR sg13g2_nor3_1
X$3045 VGND VPWR sg13g2_decap_4
X$3046 VGND ui_in[4] \$276 \$100 \$337 VPWR sg13g2_a21oi_1
X$3047 VGND ui_in[7] \$420 \$222 \$392 VPWR sg13g2_a21oi_1
X$3055 VGND ui_in[3] \$271 ui_in[0] VPWR sg13g2_nor2_1
X$3056 VGND ui_in[6] \$392 \$395 VPWR sg13g2_nor2_1
X$3057 VGND VPWR sg13g2_decap_8
X$3058 VGND VPWR sg13g2_decap_4
X$3060 VGND ui_in[2] ui_in[1] VPWR \$283 sg13g2_xnor2_1
X$3061 VGND VPWR sg13g2_decap_8
X$3062 VGND VPWR sg13g2_decap_8
X$3063 VGND VPWR sg13g2_decap_8
X$3064 VGND VPWR sg13g2_decap_8
X$3065 VGND VPWR sg13g2_decap_8
X$3066 VGND VPWR sg13g2_decap_8
X$3067 VGND VPWR sg13g2_decap_8
X$3068 VGND VPWR sg13g2_decap_8
X$3069 VGND VPWR sg13g2_decap_8
X$3070 VGND VPWR sg13g2_decap_8
X$3071 VGND VPWR sg13g2_decap_8
X$3072 VGND VPWR sg13g2_decap_8
X$3073 VGND VPWR sg13g2_decap_8
X$3074 VGND VPWR sg13g2_decap_8
X$3076 VGND VPWR sg13g2_decap_8
X$3077 VGND VPWR sg13g2_decap_8
X$3078 VGND VPWR sg13g2_decap_8
X$3079 VGND VPWR sg13g2_decap_8
X$3080 VGND VPWR sg13g2_decap_8
X$3081 VGND VPWR sg13g2_decap_8
X$3082 VGND VPWR sg13g2_decap_8
X$3083 VGND VPWR sg13g2_decap_8
X$3084 VGND VPWR sg13g2_decap_8
X$3085 VGND VPWR sg13g2_decap_8
X$3086 VGND VPWR sg13g2_decap_8
X$3087 VGND VPWR sg13g2_decap_8
X$3088 VGND VPWR sg13g2_decap_8
X$3089 VGND VPWR sg13g2_decap_8
X$3090 VGND VPWR sg13g2_decap_8
X$3091 VGND VPWR sg13g2_decap_8
X$3092 VGND VPWR sg13g2_decap_8
X$3093 VGND VPWR sg13g2_decap_8
X$3094 VGND VPWR sg13g2_decap_8
X$3095 VGND VPWR sg13g2_decap_8
X$3096 VGND VPWR sg13g2_decap_8
X$3097 VGND VPWR sg13g2_decap_8
X$3098 VGND VPWR sg13g2_decap_8
X$3100 VGND VPWR sg13g2_decap_4
X$3104 VGND ui_in[3] \$434 \$305 VPWR sg13g2_nor2b_1
X$3112 VGND \$435 ui_in[3] \$305 \$414 VPWR sg13g2_o21ai_1
X$3123 VGND \$457 \$419 \$110 \$357 \$249 \$435 VPWR sg13g2_a221oi_1
X$3130 VGND VPWR sg13g2_decap_8
X$3132 VGND VPWR sg13g2_decap_8
X$3135 VGND ui_in[5] \$248 ui_in[4] VPWR sg13g2_nor2b_1
X$3140 VGND VPWR sg13g2_decap_8
X$3149 VGND VPWR sg13g2_decap_8
X$3154 VGND VPWR sg13g2_decap_8
X$3156 VGND \$441 \$382 \$420 uo_out[2] VPWR sg13g2_a21o_1
X$3167 VGND VPWR sg13g2_decap_8
X$3176 VGND VPWR sg13g2_decap_4
X$3180 VGND \$386 \$442 ui_in[6] VPWR sg13g2_nand2_1
X$3190 VGND ui_in[0] \$463 \$337 VPWR sg13g2_nor2_1
X$3194 VGND VPWR sg13g2_decap_8
X$3198 VGND VPWR sg13g2_decap_8
X$3201 VGND \$446 \$52 \$65 \$465 VPWR sg13g2_a21o_1
X$3204 VGND VPWR sg13g2_decap_8
X$3210 VGND VPWR sg13g2_decap_8
X$3221 VGND VPWR sg13g2_decap_8
X$3231 VGND \$271 \$451 \$38 VPWR sg13g2_nand2_1
X$3238 VGND VPWR sg13g2_decap_4
X$3243 VGND \$395 \$452 \$424 \$271 VPWR sg13g2_nor3_1
X$3251 VGND \$283 \$424 ui_in[3] VPWR sg13g2_nor2b_1
X$3253 VGND VPWR sg13g2_decap_8
X$3259 VGND ui_in[3] \$337 ui_in[1] VPWR sg13g2_and2_1
X$3267 VGND VPWR sg13g2_decap_8
X$3268 VGND VPWR sg13g2_decap_8
X$3269 VGND VPWR sg13g2_decap_8
X$3270 VGND VPWR sg13g2_decap_8
X$3271 VGND VPWR sg13g2_decap_8
X$3272 VGND VPWR sg13g2_decap_8
X$3273 VGND VPWR sg13g2_decap_8
X$3274 VGND VPWR sg13g2_decap_8
X$3276 VGND VPWR sg13g2_decap_8
X$3277 VGND VPWR sg13g2_decap_8
X$3278 VGND VPWR sg13g2_decap_8
X$3279 VGND VPWR sg13g2_decap_8
X$3280 VGND VPWR sg13g2_decap_8
X$3281 VGND VPWR sg13g2_decap_8
X$3285 VGND VPWR sg13g2_decap_8
X$3286 VGND VPWR sg13g2_decap_8
X$3287 VGND VPWR sg13g2_decap_8
X$3288 VGND VPWR sg13g2_decap_8
X$3289 VGND VPWR sg13g2_decap_8
X$3290 VGND VPWR sg13g2_decap_8
X$3291 VGND VPWR sg13g2_decap_8
X$3292 VGND VPWR sg13g2_decap_8
X$3293 VGND VPWR sg13g2_decap_8
X$3294 VGND VPWR sg13g2_decap_8
X$3295 VGND VPWR sg13g2_decap_8
X$3296 VGND VPWR sg13g2_decap_8
X$3297 VGND VPWR sg13g2_decap_8
X$3298 VGND VPWR sg13g2_decap_8
X$3299 VGND VPWR sg13g2_decap_8
X$3300 VGND VPWR sg13g2_decap_8
X$3301 VGND VPWR sg13g2_decap_8
X$3302 VGND VPWR sg13g2_decap_8
X$3303 VGND VPWR sg13g2_decap_8
X$3304 VGND VPWR sg13g2_decap_8
X$3305 VGND VPWR sg13g2_decap_8
X$3306 VGND VPWR sg13g2_decap_8
X$3307 VGND VPWR sg13g2_decap_8
X$3311 VGND VPWR sg13g2_decap_8
X$3320 VGND \$305 \$549 ui_in[3] VPWR sg13g2_nand2b_1
X$3324 VGND VPWR sg13g2_decap_4
X$3330 VGND \$519 ui_in[6] \$249 \$549 ui_in[5] \$111 VPWR sg13g2_a221oi_1
X$3339 VGND \$457 \$467 ui_in[7] VPWR sg13g2_or2_1
X$3340 VGND uo_out[4] \$519 \$467 \$520 VPWR sg13g2_o21ai_1
X$3342 VGND VPWR sg13g2_decap_8
X$3350 VGND \$587 \$468 ui_in[6] \$248 \$522 VPWR sg13g2_nor4_1
X$3352 VGND \$468 \$434 \$323 \$523 VPWR sg13g2_nor3_1
X$3354 VGND ui_in[4] \$523 ui_in[5] VPWR sg13g2_or2_1
X$3357 VGND \$523 \$472 ui_in[3] ui_in[2] VPWR sg13g2_a21oi_1
X$3360 VGND ui_in[6] \$546 \$384 \$472 VPWR sg13g2_a21oi_1
X$3365 VGND \$500 \$441 \$525 VPWR sg13g2_nor2_1
X$3368 VGND ui_in[5] \$558 \$463 VPWR sg13g2_nor2_1
X$3372 VGND \$599 \$442 \$558 \$480 \$110 \$465 VPWR sg13g2_a221oi_1
X$3379 VGND \$384 ui_in[1] \$411 \$505 VPWR sg13g2_o21ai_1
X$3382 VGND ui_in[4] \$480 \$411 \$337 VPWR sg13g2_a21oi_1
X$3385 VGND \$92 \$505 ui_in[1] VPWR sg13g2_nand2_1
X$3389 VGND \$505 \$446 \$568 VPWR sg13g2_nor2b_1
X$3397 VGND \$189 \$619 \$568 \$500 VPWR sg13g2_a21oi_1
X$3400 VGND ui_in[3] \$568 \$135 VPWR sg13g2_nor2_1
X$3402 VGND \$283 \$500 \$253 VPWR sg13g2_nand2_1
X$3405 VGND ui_in[5] \$484 VPWR sg13g2_inv_1
X$3406 VGND \$522 \$484 \$271 \$283 \$100 \$337 VPWR sg13g2_a221oi_1
X$3415 VGND \$495 \$484 ui_in[4] \$489 \$480 \$451 VPWR sg13g2_a221oi_1
X$3417 VGND VPWR sg13g2_decap_8
X$3433 VGND ui_in[4] \$100 \$337 \$491 VPWR sg13g2_a21o_1
X$3435 VGND \$274 \$283 \$492 \$253 \$489 VPWR sg13g2_a22oi_1
X$3442 VGND ui_in[3] \$492 ui_in[0] VPWR sg13g2_nor2b_1
X$3443 VGND VPWR sg13g2_decap_8
X$3444 VGND VPWR sg13g2_decap_8
X$3445 VGND VPWR sg13g2_decap_8
X$3446 VGND VPWR sg13g2_decap_8
X$3447 VGND VPWR sg13g2_decap_8
X$3448 VGND VPWR sg13g2_decap_8
X$3449 VGND VPWR sg13g2_decap_8
X$3613 VGND VPWR sg13g2_decap_8
X$3614 VGND VPWR sg13g2_decap_8
X$3615 VGND VPWR sg13g2_decap_8
X$3616 VGND VPWR sg13g2_decap_8
X$3617 VGND VPWR sg13g2_decap_8
X$3618 VGND VPWR sg13g2_decap_8
X$3623 VGND VPWR sg13g2_decap_8
X$3624 VGND VPWR sg13g2_decap_8
X$3625 VGND VPWR sg13g2_decap_8
X$3626 VGND VPWR sg13g2_decap_8
X$3627 VGND VPWR sg13g2_decap_8
X$3628 VGND VPWR sg13g2_decap_8
X$3629 VGND VPWR sg13g2_decap_8
X$3630 VGND VPWR sg13g2_decap_8
X$3631 VGND VPWR sg13g2_decap_8
X$3632 VGND VPWR sg13g2_decap_8
X$3633 VGND VPWR sg13g2_decap_8
X$3634 VGND VPWR sg13g2_decap_8
X$3635 VGND VPWR sg13g2_decap_8
X$3636 VGND VPWR sg13g2_decap_8
X$3637 VGND VPWR sg13g2_decap_8
X$3638 VGND VPWR sg13g2_decap_8
X$3639 VGND VPWR sg13g2_decap_8
X$3640 VGND VPWR sg13g2_decap_8
X$3641 VGND VPWR sg13g2_decap_8
X$3642 VGND VPWR sg13g2_decap_8
X$3643 VGND VPWR sg13g2_decap_8
X$3644 VGND VPWR sg13g2_decap_8
X$3645 VGND VPWR sg13g2_decap_8
X$3650 VGND VPWR sg13g2_decap_4
X$3652 VGND ui_in[1] \$306 ui_in[0] VPWR sg13g2_nand2b_1
X$3654 VGND VPWR sg13g2_decap_8
X$3658 VGND VPWR sg13g2_decap_8
X$3661 VGND VPWR sg13g2_decap_4
X$3664 VGND \$525 ui_in[0] \$52 \$520 VPWR sg13g2_a21o_1
X$3668 VGND VPWR sg13g2_decap_8
X$3670 VGND VPWR sg13g2_decap_8
X$3674 VGND \$647 \$306 \$92 \$630 VPWR sg13g2_nand3_1
X$3676 VGND VPWR sg13g2_decap_4
X$3680 VGND uo_out[0] \$599 \$632 \$630 VPWR sg13g2_o21ai_1
X$3688 VGND VPWR sg13g2_decap_8
X$3692 VGND VPWR sg13g2_decap_8
X$3698 VGND \$411 \$671 \$38 \$271 VPWR sg13g2_a21oi_1
X$3708 VGND ui_in[5] \$698 \$274 \$411 VPWR sg13g2_a21oi_1
X$3717 VGND VPWR sg13g2_decap_8
X$3726 VGND VPWR sg13g2_decap_4
X$3731 VGND ui_in[7] \$632 \$634 VPWR sg13g2_nand2b_1
X$3734 VGND VPWR sg13g2_decap_4
X$3738 VGND \$634 \$619 \$569 \$661 VPWR sg13g2_o21ai_1
X$3740 VGND VPWR sg13g2_decap_8
X$3744 VGND VPWR sg13g2_decap_8
X$3751 VGND ui_in[2] \$682 ui_in[3] VPWR sg13g2_or2_1
X$3755 VGND VPWR sg13g2_decap_8
X$3756 VGND VPWR sg13g2_decap_8
X$3763 VGND \$569 \$491 \$640 ui_in[5] VPWR sg13g2_o21ai_1
X$3766 VGND \$640 \$135 \$575 ui_in[3] VPWR sg13g2_nor3_1
X$3773 VGND VPWR sg13g2_decap_8
X$3774 VGND VPWR sg13g2_decap_8
X$3775 VGND VPWR sg13g2_decap_8
X$3776 VGND VPWR sg13g2_decap_8
X$3777 VGND VPWR sg13g2_decap_8
X$3778 VGND VPWR sg13g2_decap_8
X$3779 VGND VPWR sg13g2_decap_8
X$3780 VGND VPWR sg13g2_decap_8
X$3781 VGND VPWR sg13g2_decap_4
X$3783 VGND VPWR sg13g2_decap_8
X$3784 VGND VPWR sg13g2_decap_8
X$3785 VGND VPWR sg13g2_decap_8
X$3786 VGND VPWR sg13g2_decap_8
X$3787 VGND VPWR sg13g2_decap_8
X$3788 VGND VPWR sg13g2_decap_8
X$3789 VGND VPWR sg13g2_decap_8
X$3790 VGND VPWR sg13g2_decap_8
X$3791 VGND VPWR sg13g2_decap_8
X$3792 VGND VPWR sg13g2_decap_8
X$3793 VGND VPWR sg13g2_decap_8
X$3794 VGND VPWR sg13g2_decap_8
X$3795 VGND VPWR sg13g2_decap_8
X$3796 VGND VPWR sg13g2_decap_8
X$3797 VGND VPWR sg13g2_decap_8
X$3798 VGND VPWR sg13g2_decap_8
X$3799 VGND VPWR sg13g2_decap_8
X$3800 VGND VPWR sg13g2_decap_8
X$3801 VGND VPWR sg13g2_decap_8
X$3802 VGND VPWR sg13g2_decap_8
X$3803 VGND VPWR sg13g2_decap_8
X$3804 VGND VPWR sg13g2_decap_8
X$3805 VGND VPWR sg13g2_decap_8
X$3806 VGND VPWR sg13g2_decap_8
X$3807 VGND VPWR sg13g2_decap_8
X$3808 VGND VPWR sg13g2_decap_8
X$3809 VGND VPWR sg13g2_decap_8
X$3810 VGND VPWR sg13g2_decap_8
X$3811 VGND VPWR sg13g2_decap_8
X$3813 VGND ui_in[0] \$707 ui_in[1] VPWR sg13g2_nor2b_1
X$3815 VGND uo_out[7] \$38 \$525 \$707 VPWR sg13g2_nor3_1
X$3819 VGND \$750 \$100 \$707 \$647 VPWR sg13g2_o21ai_1
X$3822 VGND ui_in[6] \$647 \$710 VPWR sg13g2_and2_1
X$3823 VGND \$710 \$525 ui_in[6] VPWR sg13g2_nand2_1
X$3824 VGND VPWR sg13g2_decap_4
X$3828 VGND \$647 \$253 ui_in[1] \$665 VPWR sg13g2_nand3_1
X$3832 VGND \$227 uo_out[3] \$665 VPWR sg13g2_nand2b_1
X$3834 VGND \$44 \$716 ui_in[1] ui_in[0] VPWR sg13g2_a21oi_1
X$3835 VGND \$716 \$781 \$647 VPWR sg13g2_nand2b_1
X$3837 VGND VPWR sg13g2_decap_8
X$3844 VGND \$753 ui_in[7] \$546 \$718 \$354 \$669 VPWR sg13g2_a221oi_1
X$3849 VGND VPWR sg13g2_decap_8
X$3851 VGND ui_in[4] \$274 \$806 VPWR sg13g2_xor2_1
X$3857 VGND \$723 \$52 ui_in[3] ui_in[4] \$411 VPWR sg13g2_nor4_1
X$3862 VGND \$799 \$698 \$296 \$249 \$723 VPWR sg13g2_nor4_1
X$3865 VGND VPWR sg13g2_decap_8
X$3868 VGND ui_in[6] \$296 VPWR sg13g2_inv_1
X$3870 VGND \$677 \$777 \$249 VPWR sg13g2_or2_1
X$3874 VGND \$669 \$296 \$306 \$777 \$771 \$727 VPWR sg13g2_a221oi_1
X$3880 VGND \$688 \$729 \$410 ui_in[7] VPWR sg13g2_nor3_1
X$3881 VGND ui_in[6] \$661 \$771 \$727 VPWR sg13g2_a21oi_1
X$3886 VGND \$729 \$495 \$732 ui_in[6] VPWR sg13g2_nor3_1
X$3890 VGND \$682 \$727 \$249 VPWR sg13g2_and2_1
X$3894 VGND \$682 \$732 \$452 VPWR sg13g2_nor2b_1
X$3897 VGND \$452 \$736 \$575 \$249 VPWR sg13g2_o21ai_1
X$3901 VGND \$736 \$771 \$575 VPWR sg13g2_nand2b_1
X$3908 VGND ui_in[2] \$575 ui_in[1] VPWR sg13g2_nor2b_1
X$3912 VGND VPWR sg13g2_decap_8
X$3913 VGND VPWR sg13g2_decap_8
X$3914 VGND VPWR sg13g2_decap_8
X$3915 VGND VPWR sg13g2_decap_8
X$3916 VGND VPWR sg13g2_decap_8
X$3917 VGND VPWR sg13g2_decap_8
X$3918 VGND VPWR sg13g2_decap_8
X$3919 VGND VPWR sg13g2_decap_8
X$4087 VGND VPWR sg13g2_decap_8
X$4088 VGND VPWR sg13g2_decap_8
X$4089 VGND VPWR sg13g2_decap_8
X$4090 VGND VPWR sg13g2_decap_8
X$4091 VGND VPWR sg13g2_decap_8
X$4092 VGND VPWR sg13g2_decap_8
X$4094 VGND VPWR sg13g2_decap_8
X$4095 VGND VPWR sg13g2_decap_8
X$4096 VGND VPWR sg13g2_decap_8
X$4097 VGND VPWR sg13g2_decap_8
X$4098 VGND VPWR sg13g2_decap_8
X$4101 VGND uio_oe[7] \$779 VPWR sg13g2_buf_1
X$4102 VGND uio_oe[6] \$779 VPWR sg13g2_buf_1
X$4103 VGND \$779 VPWR sg13g2_tielo
X$4105 VGND uio_oe[5] \$779 VPWR sg13g2_buf_1
X$4106 VGND VPWR sg13g2_decap_4
X$4107 VGND uio_oe[4] \$779 VPWR sg13g2_buf_1
X$4108 VGND VPWR sg13g2_decap_4
X$4109 VGND uio_oe[3] \$779 VPWR sg13g2_buf_1
X$4110 VGND VPWR sg13g2_decap_4
X$4111 VGND uio_oe[2] \$779 VPWR sg13g2_buf_1
X$4114 VGND uio_oe[1] \$779 VPWR sg13g2_buf_1
X$4115 VGND VPWR sg13g2_decap_4
X$4116 VGND uio_oe[0] \$779 VPWR sg13g2_buf_1
X$4117 VGND VPWR sg13g2_decap_4
X$4118 VGND uio_out[7] \$779 VPWR sg13g2_buf_1
X$4119 VGND VPWR sg13g2_decap_4
X$4121 VGND uio_out[6] \$779 VPWR sg13g2_buf_1
X$4122 VGND VPWR sg13g2_decap_4
X$4123 VGND uio_out[5] \$779 VPWR sg13g2_buf_1
X$4124 VGND VPWR sg13g2_decap_4
X$4125 VGND uio_out[4] \$779 VPWR sg13g2_buf_1
X$4128 VGND uio_out[3] \$779 VPWR sg13g2_buf_1
X$4129 VGND VPWR sg13g2_decap_4
X$4130 VGND uio_out[2] \$779 VPWR sg13g2_buf_1
X$4131 VGND VPWR sg13g2_decap_4
X$4132 VGND uio_out[1] \$779 VPWR sg13g2_buf_1
X$4133 VGND uio_out[0] \$779 VPWR sg13g2_buf_1
X$4134 VGND VPWR sg13g2_decap_8
X$4136 VGND VPWR sg13g2_decap_8
X$4137 VGND VPWR sg13g2_decap_4
X$4138 VGND \$753 uo_out[6] \$750 VPWR sg13g2_nand2b_1
X$4143 VGND ui_in[7] ui_in[5] ui_in[3] \$710 ui_in[4] VPWR sg13g2_and4_1
X$4145 VGND VPWR sg13g2_decap_8
X$4146 VGND VPWR sg13g2_decap_8
X$4151 VGND VPWR sg13g2_decap_4
X$4153 VGND uo_out[5] \$587 \$802 \$781 VPWR sg13g2_o21ai_1
X$4158 VGND \$688 uo_out[1] uo_out[7] VPWR sg13g2_or2_1
X$4160 VGND VPWR sg13g2_decap_4
X$4162 VGND \$799 \$802 ui_in[7] VPWR sg13g2_or2_1
X$4164 VGND VPWR sg13g2_decap_8
X$4165 VGND VPWR sg13g2_decap_8
X$4166 VGND \$718 \$671 \$806 ui_in[5] VPWR sg13g2_o21ai_1
X$4168 VGND VPWR sg13g2_decap_4
X$4169 VGND ui_in[2] \$411 ui_in[0] VPWR sg13g2_and2_1
X$4170 VGND VPWR sg13g2_decap_8
X$4173 VGND VPWR sg13g2_decap_8
X$4175 VGND VPWR sg13g2_decap_8
X$4177 VGND \$677 ui_in[1] ui_in[4] ui_in[3] VPWR sg13g2_nor3_1
X$4179 VGND VPWR sg13g2_decap_8
X$4180 VGND VPWR sg13g2_decap_8
X$4182 VGND VPWR sg13g2_decap_8
X$4184 VGND VPWR sg13g2_decap_8
X$4187 VGND VPWR sg13g2_decap_4
X$4189 VGND ui_in[5] \$249 ui_in[4] VPWR sg13g2_nor2_1
X$4190 VGND ui_in[0] \$736 ui_in[3] VPWR sg13g2_nand2_1
X$4191 VGND ui_in[3] \$274 ui_in[1] VPWR sg13g2_nor2_1
X$4193 VGND VPWR sg13g2_decap_8
X$4194 VGND VPWR sg13g2_decap_8
X$4195 VGND VPWR sg13g2_decap_8
X$4196 VGND VPWR sg13g2_decap_8
X$4197 VGND VPWR sg13g2_decap_8
X$4198 VGND VPWR sg13g2_decap_8
X$4199 VGND VPWR sg13g2_decap_8
X$4200 VGND VPWR sg13g2_decap_8
X$4201 VGND VPWR sg13g2_decap_4
.ENDS tt_um_chip_rom

.SUBCKT sg13g2_tielo VSS L_LO VDD
XM$1 VSS \$6 \$5 VSS sg13_lv_nmos L=0.13u W=0.385u AS=0.305425p AD=0.1309p
+ PS=2.07u PD=1.45u
XM$2 VSS \$3 L_LO VSS sg13_lv_nmos L=0.13u W=0.88u AS=0.305425p AD=0.2992p
+ PS=2.07u PD=2.44u
XM$3 VDD \$6 \$6 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.326925p AD=0.102p
+ PS=2.255u PD=1.28u
XM$4 VDD \$5 \$3 VDD sg13_lv_pmos L=0.13u W=1.045u AS=0.326925p AD=0.3553p
+ PS=2.255u PD=2.77u
.ENDS sg13g2_tielo

.SUBCKT sg13g2_buf_1 VSS \$2 \$3 VDD
XM$1 VSS \$3 \$4 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.159375p AD=0.247625p
+ PS=1.19u PD=2.29u
XM$2 VSS \$4 \$2 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.159375p AD=0.2516p
+ PS=1.19u PD=2.16u
XM$3 VDD \$3 \$4 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2051p AD=0.3024p PS=1.52u
+ PD=2.4u
XM$4 VDD \$4 \$2 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2051p AD=0.4032p PS=1.52u
+ PD=2.96u
.ENDS sg13g2_buf_1

.SUBCKT sg13g2_or3_1 VSS C B A X VDD
XM$1 \$3 C VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.187p AD=0.1045p PS=1.78u
+ PD=0.93u
XM$2 VSS B \$3 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.1045p AD=0.198p PS=0.93u
+ PD=1.27u
XM$3 \$3 A VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.198p AD=0.13395p PS=1.27u
+ PD=1.12u
XM$4 VSS \$3 X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.13395p AD=0.2516p PS=1.12u
+ PD=2.16u
XM$5 \$3 C \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.1275p PS=2.68u
+ PD=1.255u
XM$6 \$9 B \$8 VDD sg13_lv_pmos L=0.13u W=1u AS=0.1275p AD=0.22p PS=1.255u
+ PD=1.44u
XM$7 \$8 A VDD VDD sg13_lv_pmos L=0.13u W=1u AS=0.22p AD=0.3822p PS=1.44u
+ PD=1.84u
XM$8 VDD \$3 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3822p AD=0.3808p PS=1.84u
+ PD=2.92u
.ENDS sg13g2_or3_1

.SUBCKT sg13g2_and4_1 VSS A B C X D VDD
XM$1 \$2 A \$9 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p AD=0.0832p PS=1.96u
+ PD=0.9u
XM$2 \$9 B \$8 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.0832p AD=0.0832p PS=0.9u
+ PD=0.9u
XM$3 \$8 C \$10 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.0832p AD=0.1408p PS=0.9u
+ PD=1.08u
XM$4 \$10 D VSS VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1408p AD=0.1351p PS=1.08u
+ PD=1.12u
XM$5 VSS \$2 X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1351p AD=0.3552p PS=1.12u
+ PD=2.44u
XM$6 VDD A \$2 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p AD=0.1596p PS=2.36u
+ PD=1.22u
XM$7 \$2 B VDD VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1596p AD=0.1596p PS=1.22u
+ PD=1.22u
XM$8 VDD C \$2 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1596p AD=0.1848p PS=1.22u
+ PD=1.28u
XM$9 VDD D \$2 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2044p AD=0.1848p PS=1.53u
+ PD=1.28u
XM$10 VDD \$2 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2044p AD=0.5376p PS=1.53u
+ PD=3.2u
.ENDS sg13g2_and4_1

.SUBCKT sg13g2_nor4_1 VSS Y C A B D VDD
XM$1 VSS A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u
+ PD=1.12u
XM$2 Y B VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.1406p PS=1.12u
+ PD=1.12u
XM$3 VSS C Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.1406p PS=1.12u
+ PD=1.12u
XM$4 Y D VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.237575p PS=1.12u
+ PD=2.16u
XM$5 VDD A \$8 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.1624p PS=2.92u
+ PD=1.41u
XM$6 \$8 B \$9 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1624p AD=0.2464p PS=1.41u
+ PD=1.56u
XM$7 \$9 C \$10 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2464p AD=0.2464p PS=1.56u
+ PD=1.56u
XM$8 \$10 D Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2464p AD=0.4032p PS=1.56u
+ PD=2.96u
.ENDS sg13g2_nor4_1

.SUBCKT sg13g2_nand3b_1 VSS A_N C Y B VDD
XM$1 VSS A_N \$2 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.1839p AD=0.187p PS=1.255u
+ PD=1.78u
XM$2 VSS C \$8 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1839p AD=0.1739p PS=1.255u
+ PD=1.21u
XM$3 \$8 B \$7 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1739p AD=0.10915p PS=1.21u
+ PD=1.035u
XM$4 \$7 \$2 Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.10915p AD=0.3404p PS=1.035u
+ PD=2.4u
XM$5 \$2 A_N VDD VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p AD=0.2198p PS=2.36u
+ PD=1.53u
XM$6 VDD C Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2198p AD=0.2128p PS=1.53u
+ PD=1.5u
XM$7 Y B VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u
+ PD=1.5u
XM$8 VDD \$2 Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_nand3b_1

.SUBCKT sg13g2_xnor2_1 VSS A B VDD Y
XM$1 VSS A \$6 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2272p AD=0.0784p PS=1.99u
+ PD=0.885u
XM$2 \$6 B \$3 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.0784p AD=0.2176p PS=0.885u
+ PD=1.96u
XM$3 VSS A \$5 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1898p AD=0.2516p PS=1.36u
+ PD=2.16u
XM$4 VSS B \$5 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1898p AD=0.1406p PS=1.36u
+ PD=1.12u
XM$5 \$5 \$3 Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u
+ PD=2.16u
XM$6 VDD A \$3 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.4536p AD=0.1596p PS=2.76u
+ PD=1.22u
XM$7 VDD B \$3 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2891p AD=0.1596p PS=1.695u
+ PD=1.22u
XM$8 VDD A \$9 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2891p AD=0.1428p PS=1.695u
+ PD=1.375u
XM$9 \$9 B Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1428p AD=0.2408p PS=1.375u
+ PD=1.55u
XM$10 Y \$3 VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2408p AD=0.3808p PS=1.55u
+ PD=2.92u
.ENDS sg13g2_xnor2_1

.SUBCKT sg13g2_a21o_1 VSS B1 A1 A2 X VDD
XM$1 X \$2 VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2351p AD=0.15745p PS=2.16u
+ PD=1.175u
XM$2 VSS B1 \$2 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.15745p AD=0.1216p
+ PS=1.175u PD=1.02u
XM$3 \$2 A1 \$7 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1216p AD=0.0816p PS=1.02u
+ PD=0.895u
XM$4 \$7 A2 VSS VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.0816p AD=0.2176p PS=0.895u
+ PD=1.96u
XM$5 \$2 B1 \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.35p AD=0.2125p PS=2.7u
+ PD=1.425u
XM$6 \$9 A1 VDD VDD sg13_lv_pmos L=0.13u W=1u AS=0.2125p AD=0.19p PS=1.425u
+ PD=1.38u
XM$7 VDD A2 \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.19p AD=0.34p PS=1.38u PD=2.68u
XM$8 X \$2 VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.3808p PS=2.92u
+ PD=2.92u
.ENDS sg13g2_a21o_1

.SUBCKT sg13g2_a22oi_1 VSS A1 B1 B2 A2 Y VDD
XM$1 VSS B1 \$8 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2553p AD=0.13875p PS=2.17u
+ PD=1.115u
XM$2 \$8 B2 Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.13875p AD=0.2664p PS=1.115u
+ PD=1.46u
XM$3 Y A1 \$7 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2664p AD=0.0962p PS=1.46u
+ PD=1u
XM$4 \$7 A2 VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.0962p AD=0.2516p PS=1u
+ PD=2.16u
XM$5 VDD A1 \$10 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2716p PS=2.92u
+ PD=1.605u
XM$6 \$10 B1 Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2716p AD=0.2128p PS=1.605u
+ PD=1.5u
XM$7 Y B2 \$10 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2744p PS=1.5u
+ PD=1.61u
XM$8 \$10 A2 VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2744p AD=0.3808p PS=1.61u
+ PD=2.92u
.ENDS sg13g2_a22oi_1

.SUBCKT sg13g2_inv_1 VSS A Y VDD
XM$1 VSS A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p AD=0.259p PS=2.18u
+ PD=2.18u
XM$2 VDD A Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p AD=0.392p PS=2.94u
+ PD=2.94u
.ENDS sg13g2_inv_1

.SUBCKT sg13g2_or2_1 VSS B X A VDD
XM$1 VSS B \$4 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.187p AD=0.1045p PS=1.78u
+ PD=0.93u
XM$2 \$4 A VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.1045p AD=0.1469p PS=0.93u
+ PD=1.155u
XM$3 VSS \$4 X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1469p AD=0.2516p PS=1.155u
+ PD=2.16u
XM$4 \$4 B \$7 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p AD=0.1596p PS=2.36u
+ PD=1.22u
XM$5 VDD A \$7 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2226p AD=0.1596p PS=1.535u
+ PD=1.22u
XM$6 VDD \$4 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2226p AD=0.3976p PS=1.535u
+ PD=2.95u
.ENDS sg13g2_or2_1

.SUBCKT sg13g2_and2_1 VSS A X B VDD
XM$1 \$3 A \$6 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p AD=0.1216p PS=1.96u
+ PD=1.02u
XM$2 VSS B \$6 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p AD=0.1216p PS=1.12u
+ PD=1.02u
XM$3 VSS \$3 X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1331p AD=0.2516p PS=1.12u
+ PD=2.16u
XM$4 VDD A \$3 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p AD=0.1596p PS=2.36u
+ PD=1.22u
XM$5 VDD B \$3 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p AD=0.1596p PS=1.5u
+ PD=1.22u
XM$6 VDD \$3 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1918p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_and2_1

.SUBCKT sg13g2_nor2b_1 VSS B_N Y A VDD
XM$1 VSS B_N \$5 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.17255p AD=0.187p PS=1.25u
+ PD=1.78u
XM$2 VSS \$5 Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.17255p AD=0.1406p PS=1.25u
+ PD=1.12u
XM$3 Y A VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u
+ PD=2.16u
XM$4 \$5 B_N VDD VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p AD=0.2618p PS=2.36u
+ PD=1.63u
XM$5 VDD \$5 \$7 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2618p AD=0.1176p PS=1.63u
+ PD=1.33u
XM$6 \$7 A Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p AD=0.3808p PS=1.33u
+ PD=2.92u
.ENDS sg13g2_nor2b_1

.SUBCKT sg13g2_a221oi_1 \$1 \$2 \$3 \$4 \$5 \$6 \$7 \$10
XM$1 \$2 \$6 \$9 \$1 sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u
+ PD=1.12u
XM$2 \$9 \$7 \$1 \$1 sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u
+ PD=2.16u
XM$3 \$2 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u
+ PD=1.12u
XM$4 \$1 \$4 \$8 \$1 sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.1406p PS=1.12u
+ PD=1.12u
XM$5 \$8 \$5 \$2 \$1 sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u
+ PD=2.16u
XM$6 \$10 \$6 \$12 \$10 sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p
+ PS=2.92u PD=1.5u
XM$7 \$12 \$7 \$10 \$10 sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p
+ PS=1.5u PD=2.92u
XM$8 \$2 \$3 \$11 \$10 sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p
+ PS=2.92u PD=1.5u
XM$9 \$11 \$4 \$12 \$10 sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p
+ PS=1.5u PD=1.5u
XM$10 \$12 \$5 \$11 \$10 sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p
+ PS=1.5u PD=2.92u
.ENDS sg13g2_a221oi_1

.SUBCKT sg13g2_decap_4 VSS VDD
XM$1 VSS VDD VSS VSS sg13_lv_nmos L=1u W=0.42u AS=0.1428p AD=0.1428p PS=1.52u
+ PD=1.52u
XM$2 VDD VSS VDD VDD sg13_lv_pmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
.ENDS sg13g2_decap_4

.SUBCKT sg13g2_nor2_1 VSS A Y B VDD
XM$1 VSS A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u
+ PD=1.12u
XM$2 Y B VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u
+ PD=2.16u
XM$3 VDD A \$6 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.4032p AD=0.1176p PS=2.96u
+ PD=1.33u
XM$4 \$6 B Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p AD=0.3808p PS=1.33u
+ PD=2.92u
.ENDS sg13g2_nor2_1

.SUBCKT sg13g2_nor3_1 VSS Y B C A VDD
XM$1 VSS A Y VSS sg13_lv_nmos L=0.13u W=0.77u AS=0.2618p AD=0.1694p PS=2.22u
+ PD=1.21u
XM$2 Y B VSS VSS sg13_lv_nmos L=0.13u W=0.77u AS=0.1694p AD=0.1463p PS=1.21u
+ PD=1.15u
XM$3 VSS C Y VSS sg13_lv_nmos L=0.13u W=0.77u AS=0.1463p AD=0.2618p PS=1.15u
+ PD=2.22u
XM$4 VDD A \$7 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.1764p PS=2.92u
+ PD=1.435u
XM$5 \$7 B \$8 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1764p AD=0.182p PS=1.435u
+ PD=1.445u
XM$6 \$8 C Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.182p AD=0.3808p PS=1.445u
+ PD=2.92u
.ENDS sg13g2_nor3_1

.SUBCKT sg13g2_nand2_1 VSS B Y A VDD
XM$1 VSS B \$5 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.0666p PS=2.16u
+ PD=0.92u
XM$2 \$5 A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.0666p AD=0.2516p PS=0.92u
+ PD=2.16u
XM$3 VDD B Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
XM$4 Y A VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_nand2_1

.SUBCKT sg13g2_a21oi_1 VSS B1 Y A1 A2 VDD
XM$1 VSS B1 Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u
+ PD=1.12u
XM$2 Y A1 \$6 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.1406p PS=1.12u
+ PD=1.12u
XM$3 \$6 A2 VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u
+ PD=2.16u
XM$4 Y B1 \$8 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
XM$5 \$8 A1 VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u
+ PD=1.5u
XM$6 VDD A2 \$8 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_a21oi_1

.SUBCKT sg13g2_decap_8 VSS VDD
XM$1 VSS VDD VSS VSS sg13_lv_nmos L=1u W=0.84u AS=0.2226p AD=0.2226p PS=2.32u
+ PD=2.32u
XM$3 VDD VSS VDD VDD sg13_lv_pmos L=1u W=2u AS=0.53p AD=0.53p PS=4.06u PD=4.06u
.ENDS sg13g2_decap_8

.SUBCKT sg13g2_nand2b_1 VSS A_N Y B VDD
XM$1 VSS A_N \$3 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.25975p AD=0.187p PS=1.46u
+ PD=1.78u
XM$2 VSS B \$6 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.25975p AD=0.0666p PS=1.46u
+ PD=0.92u
XM$3 \$6 \$3 Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.0666p AD=0.2516p PS=0.92u
+ PD=2.16u
XM$4 \$3 A_N VDD VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p AD=0.2198p PS=2.36u
+ PD=1.53u
XM$5 VDD B Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2198p AD=0.2128p PS=1.53u
+ PD=1.5u
XM$6 Y \$3 VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_nand2b_1

.SUBCKT sg13g2_nand3_1 VSS C B A Y VDD
XM$1 VSS C \$6 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2886p AD=0.17205p PS=2.26u
+ PD=1.205u
XM$2 \$6 B \$7 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.17205p AD=0.10915p
+ PS=1.205u PD=1.035u
XM$3 \$7 A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.10915p AD=0.3293p PS=1.035u
+ PD=2.37u
XM$4 VDD C Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
XM$5 Y B VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u
+ PD=1.5u
XM$6 VDD A Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_nand3_1

.SUBCKT sg13g2_nand4_1 VSS D C B A VDD Y
XM$1 VSS D \$8 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2886p AD=0.13875p PS=2.26u
+ PD=1.115u
XM$2 \$8 C \$7 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.13875p AD=0.14245p
+ PS=1.115u PD=1.125u
XM$3 \$7 B \$6 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.14245p AD=0.1406p PS=1.125u
+ PD=1.12u
XM$4 \$6 A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u
+ PD=2.16u
XM$5 VDD D Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
XM$6 Y C VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u
+ PD=1.5u
XM$7 VDD B Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u
+ PD=1.5u
XM$8 Y A VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_nand4_1

.SUBCKT sg13g2_o21ai_1 VSS Y A1 A2 B1 VDD
XM$1 \$2 A1 VSS VSS sg13_lv_nmos L=0.15u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u
+ PD=1.12u
XM$2 VSS A2 \$2 VSS sg13_lv_nmos L=0.15u W=0.74u AS=0.1406p AD=0.1406p PS=1.12u
+ PD=1.12u
XM$3 \$2 B1 Y VSS sg13_lv_nmos L=0.15u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u
+ PD=2.16u
XM$4 VDD A1 \$8 VDD sg13_lv_pmos L=0.15u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
XM$5 \$8 A2 Y VDD sg13_lv_pmos L=0.15u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u
+ PD=1.5u
XM$6 Y B1 VDD VDD sg13_lv_pmos L=0.15u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_o21ai_1

.SUBCKT sg13g2_xor2_1 VSS A B X VDD
XM$1 VSS A \$5 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.374p AD=0.174625p PS=2.46u
+ PD=1.185u
XM$2 VSS B \$5 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.15245p AD=0.174625p
+ PS=1.17u PD=1.185u
XM$3 VSS A \$6 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.15245p AD=0.0888p PS=1.17u
+ PD=0.98u
XM$4 \$6 B X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.0888p AD=0.1628p PS=0.98u
+ PD=1.18u
XM$5 X \$5 VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1628p AD=0.3108p PS=1.18u
+ PD=2.32u
XM$6 \$8 A VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
XM$7 VDD B \$8 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u
+ PD=1.5u
XM$8 \$8 \$5 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
XM$9 VDD A \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.36p AD=0.1225p PS=2.72u
+ PD=1.245u
XM$10 \$9 B \$5 VDD sg13_lv_pmos L=0.13u W=1u AS=0.1225p AD=0.34p PS=1.245u
+ PD=2.68u
.ENDS sg13g2_xor2_1

* Tiny Tapeout ROM testbench
* Run with `make sim_nand`

.include "pdk_lib.spice"

* Power supply
V1 VGND 0 0
V2 VPWR VGND 1.2

.include "tt_um_chip_rom.spice"

x1 VGND VPWR clk ena rst_n
+ addr0 addr1 addr2 addr3 addr4 addr5 addr6 addr7
+ VGND VGND VGND VGND VGND VGND VGND VGND
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ data0 data1 data2 data3 data4 data5 data6 data7
+ tt_um_chip_rom

* Tie the clock to ground, ena/rst_n to power
Vtie_clk clk 0 0
Vtie_ena ena VPWR 0
Vtie_rst_n rst_n VPWR 0

* Iterate over all possible ROM addresses
V3  addr0 VGND PULSE(0 1.8 10n  0 0 10n  20n)
V4  addr1 VGND PULSE(0 1.8 20n  0 0 20n  40n)
V5  addr2 VGND PULSE(0 1.8 40n  0 0 40n  80n)
V6  addr3 VGND PULSE(0 1.8 80n  0 0 80n  160n)
V7  addr4 VGND PULSE(0 1.8 160n 0 0 160n 320n)
V8  addr5 VGND PULSE(0 1.8 320n 0 0 320n 640n)
V9  addr6 VGND PULSE(0 1.8 640n 0 0 640n 1280n)
V10 addr7 VGND PULSE(0 1.8 1280n 0 0 1280n 2560n)

.param mc_mm_switch=0

.tran 5n 2560n

.control
run
set wr_vecnames
set wr_singlescale
wrdata rom_signals.txt addr0 addr1 addr2 addr3 addr4 addr5 addr6 addr7 data0 data1 data2 data3 data4 data5 data6 data7
.endc
.end

.end
